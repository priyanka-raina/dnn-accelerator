
//------> /hd/cad/mentor/2016.9/Mgc_home/pkgs/siflibs/mgc_out_stdreg_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule



//------> /hd/cad/mentor/2016.9/Mgc_home/pkgs/siflibs/mgc_io_sync_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v1 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


module mgc_in_sync_v1 (vd, vz);
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule



//------> /hd/cad/mentor/2016.9/Mgc_home/pkgs/siflibs/mgc_in_wire_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule


//------> /hd/cad/mentor/2016.9/Mgc_home/pkgs/siflibs/designcompiler/28nm.verilog.v 
 
`ifdef __core__ 

`else 

`define __core__ 

module core (
				acc,
				addra,
				addrb,
				clamp_mem,
				clk,
				csa_n,
				csb_n,
				dinb,
				douta,
				scan_n,
				shift_n,
				sin,
				slp_nret_n,
				slp_ret_n,
				sout
			);
   // Parameter declarations
   parameter filename = "NONE";
   //parameter filename_size = 128;
   parameter SCAN_DEPTH_ADDR = 9;
   parameter WORDS = 256;
   parameter ADDR_WIDTH = 8;
   parameter BPW = 64;
   //parameter WORDX = {BPW{1'bx}};
   parameter FAILED_IO = 0;
   parameter FAILED_ADDR = 0;
   parameter ACC_DEBUG = 0;

   // Output and Input ports
   input	[3:0]	acc ;
   input	[7:0]	addra ;
   input	[7:0]	addrb ;
   input		clamp_mem ;
   input		clk ;
   input		csa_n ;
   input		csb_n ;
   input	[63:0]	dinb ;
   output	[63:0]	douta ;
   input		scan_n ;
   input		shift_n ;
   input		sin ;
   input		slp_nret_n ;
   input		slp_ret_n ;
   output		sout ;

   // Internal registers and memory array definitions
   reg                                                            prev_clk;
   reg [BPW - 1:0]                                                douta;
   reg                                                            sout;
   reg [BPW - 1:0]                                                Dinb;
   reg                                                            Csa_n;
   reg                                                            Csb_n;
   reg [BPW - 1:0]                                                Wbtb_n;
   reg [SCAN_DEPTH_ADDR :0]				          Addra;
   reg [SCAN_DEPTH_ADDR :0]				          Addrb;
   reg [SCAN_DEPTH_ADDR :0]				          Addra_r;
   reg [SCAN_DEPTH_ADDR :0]				          Addrb_r;
   reg [SCAN_DEPTH_ADDR :0]				          Addra_rw;
   reg [SCAN_DEPTH_ADDR :0]				          Addrb_rw;
   reg [BPW - 1:0]                                                Dinb_r;
   reg                                                            Csa_n_r;
   reg                                                            Csb_n_r;
   reg [BPW - 1:0]                                                Wbtb_n_r;
   reg                                                            wait_period;
   reg  	            			                  slp_min_period;
   reg                                                            flag_tpd4;
   reg                                                            flag_tpd1;
   reg [BPW - 1:0]                                                temp_write_reg;
   reg [BPW - 1:0]                                                temp_read_reg;
   reg [BPW - 1:0]                                                i_memArray [WORDS - 1:0];

   reg [BPW - 1:0]                                                wbtb_n;
   reg [2*BPW + 2*SCAN_DEPTH_ADDR + 1 : 0 ]            	  	  scan_reg;

   reg                                                            functional_mode;
   reg                                                            read_op;
   reg                                                            write_op;

   reg                                                            scan_op;

   reg                                                            dummy_clock_reg;
   reg                                                            prev_slp_nret_n;

   reg                                                            prev_clamp_mem;

   reg [8*128 - 1:0]                                    MEMORY_TRACE_LOG = "off";
   reg [8*128 - 1:0]                                    IMAGE_FILE = "NULL";
   reg                                                            NO_WARNING = 0;
   reg                                                            NO_CORRUPT = 0;
   reg                           		                  valid_acc = 0 ;
   integer                                                        log_file, image_file,count;
   reg                           		                  FAILURE_INJECT = 0 ;
   reg [BPW - 1:0] 	     	 				  temp_write_failure_reg;       // used for failure injection
   reg [5: 0]                           		          failed_io;
   reg [ADDR_WIDTH -1 : 0]                          failed_addr;
   time                                                        	prev_time, current_time, diff_time, sleep_time; 
   // Getting the memory modes
   task check_mode;
      begin
    // Adding waitperiod here to make sure nothing happens in wait period.. (dummy_clock_reg added for the same reason..) 
        functional_mode = scan_n & shift_n & dummy_clock_reg & ~clamp_mem & valid_acc & slp_ret_n & slp_nret_n;
        read_op = scan_n & shift_n & dummy_clock_reg & ~clamp_mem & valid_acc & slp_ret_n & slp_nret_n & (~Csa_n_r);
        write_op = scan_n & shift_n & dummy_clock_reg & ~clamp_mem & valid_acc  & slp_ret_n & slp_nret_n & (~Csb_n_r);
        scan_op = ~scan_n & ~clamp_mem & valid_acc & slp_ret_n & slp_nret_n;
      end
   endtask

   // Write all 1's into wbt_n for word writable memory
   task get_wbtb_for_word;
      // Loop Counter
      integer 	i;
      begin
         for (i = 0; i < BPW; i = i + 1)
             wbtb_n[i] = 1'b0;
      end
   endtask

   task get_Addra_Addrb;
      integer i;
      integer c;
      parameter last_addr = 9;
      begin
      c = 0;
      for(i = 2; i < 5; i = i+1)
      begin
      if(i == 2)
         begin
         Addra[i] = shift_n ? addra[i] : sin ;
         Addrb[i] = shift_n ? addrb[i] : scan_reg[(2*c)] ;
         c= c+1;
         end
      else if((i > 2) && (i < ADDR_WIDTH)) 
         begin
         Addra[i] = shift_n ? addra[i] : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? addrb[i] : scan_reg[(2*c)] ;
         c= c+1;
         end
      else
         begin
         Addra[i] = shift_n ? 1'b0 : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? 1'b0 : scan_reg[(2*c)] ;
         c= c+1;
         end
      end

      for(i = 8; i <= 9; i = i+1)
      begin
      if(i < ADDR_WIDTH)
         begin
         Addra[i] = shift_n ? addra[i] : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? addrb[i] : scan_reg[(2*c)] ;
         c= c+1;
         end
      else
         begin
         Addra[i] = shift_n ? 1'b0 : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? 1'b0 : scan_reg[(2*c)] ;
         c= c+1;
         end
      end

      for(i = 5; i < 8; i = i+1)
      begin
      if(i < ADDR_WIDTH)
         begin
         Addra[i] = shift_n ? addra[i] : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? addrb[i] : scan_reg[(2*c)] ;
         c= c+1;
         end
      else
         begin
         Addra[i] = shift_n ? 1'b0 : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? 1'b0 : scan_reg[(2*c)] ;
         c= c+1;
         end
      end

      for(i = 0; i < 2; i = i+1)
      begin
      if(i < ADDR_WIDTH)
         begin
         Addra[i] = shift_n ? addra[i] : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? addrb[i] : scan_reg[(2*c)] ;
         c= c+1;
         end
      else
         begin
         Addra[i] = shift_n ? 1'b0 : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? 1'b0 : scan_reg[(2*c)] ;
         c= c+1;
         end
      end
   end
   endtask

   task get_Csa_n;
      begin
    Csa_n = csa_n ;
      end
   endtask

   task get_Csb_n;
      begin
    Csb_n = csb_n ;
      end
   endtask

   // Getting Din through scan logic
   // The selection is between previous scan register( width = addr_width + 1; ie 0 to addr_width; din[0] has to choose between  scan reg[addr_width] and normal din logic.  
   task get_Wbtn_n_Dinb;
      integer i;
      integer j;
      parameter C1 = 2 * SCAN_DEPTH_ADDR + 2;
      begin
	 for (i = 0; i < BPW; i = i + 1)
	   begin
	       Wbtb_n[i] = shift_n ? wbtb_n[i] : scan_reg[C1+(2*i) -1] ;
	       Dinb[i] = shift_n ? dinb[i] : scan_reg[C1+(2*i)] ;
	   end
      end
   endtask

   // Write into specified bits alone
   task bit_wise_write;
      integer i;
      begin
      for (i = 0; i < BPW; i = i + 1)
        if (!Wbtb_n_r[i])
 	 temp_write_reg[i] = Dinb_r[i];
      end
   endtask

   // Select between BIST and normal inputs
   task input_source_select;
      begin
      get_Addra_Addrb ;
      get_Csa_n ;
      get_Csb_n ;
      get_Wbtn_n_Dinb ;
      end
   endtask

   // Register inputs
   task register_inputs;
      begin
	Dinb_r     = Dinb ; 
	Addra_r    = Addra ; 
	Addrb_r    = Addrb ; 
        Wbtb_n_r   = Wbtb_n ; 
        Csa_n_r    = Csa_n ; 
        Csb_n_r    = Csb_n ; 
      end
   endtask

   // Register read/write address
   task register_rw_addr;
     parameter MSB1 = 9;
     parameter MSB2 = 8;
       begin
	 Addra_rw    = Addra_r ; 
	 Addrb_rw    = Addrb_r ; 
      end
   endtask

   // Invalidate entire memory
   task invalidate_memory;
      integer i;
      begin
         if (NO_CORRUPT == 0)
           begin
            if (NO_WARNING == 0)
              begin
              $display(" %t : Memory instance %m:: Invalidating memory contents ", $time);
              end
	    for (i = 0; i < WORDS; i = i + 1)
	       begin
	        i_memArray[i] = {BPW{1'bx}};
	       end
      end
         else
           begin
             if (NO_WARNING == 0)
               begin
                 $display("%t : Warning on memory instance %m:: NO_CORRUPT Flag is set and hence invalid inputs wont corrupt the memory !! ", $time);
               end
          end
      end
   endtask

   // Invalidate entire memory for sleep no retention
   task invalidate_memory_always;
      integer i;
      begin
	 if (NO_CORRUPT == 0)
	   begin
	    if (NO_WARNING == 0)
	      begin
	      $display(" %t : Memory instance %m:: Invalidating memory contents ", $time);
	      end
	    for (i = 0; i < WORDS; i = i + 1)
	       begin
	        i_memArray[i] = {BPW{1'bx}};
	       end
	   end
	 else
	   begin
	     if (NO_WARNING == 0)
	       begin
		 $display("%t : Warning on memory instance %m:: NO_CORRUPT Flag is set and hence sleep no retention mode wont corrupt the memory !! ", $time);
	       end
	   end
      end
   endtask

   // Clk and slp_ret_n should be zero when the clamp_mem is asserted or de-asserted
   task clamp_violation_check;
      begin
         if ((slp_ret_n !== 1'b0) && (slp_nret_n !== 1'b0))
           begin
             if (NO_WARNING == 0)
               begin
                 $display("%t : Error on memory instance %m:: Power Collapse Violation. slp_ret_n should be low ", $time);
               end
             invalidate_memory;
          end
      end
   endtask

   // memory functional cycle 
   task mem_func;
      begin
        if(wait_period == 0)
          begin
           if ( read_op == 1 )
              read ;
           if ( write_op == 1 )
              write ;
           if ((Csa_n_r === 1'bx) && ( functional_mode == 1 ))
              invalid_Csa_n_r ;
           if ((Csb_n_r === 1'bx) && ( functional_mode == 1 ))
              invalid_Csb_n_r ;
          end
      end
   endtask

   // Updating the scan chain
   task update_scan_reg;
     integer i ;
     integer j ;
     parameter C1 = 2*SCAN_DEPTH_ADDR + 2 ;
     begin
        if (scan_op == 1)
        begin
	    for (i = 0; i <= SCAN_DEPTH_ADDR; i = i + 1)
            begin
              if (i < 3)
                begin
                j = 2+i;
                scan_reg[2*i] = Addra_r[j];
                scan_reg[(2*i)+1] = Addrb_r[j];
                end
              else if ((i == 3) || (i == 4))
                begin
                j = 9-4+i;
                scan_reg[2*i] = Addra_r[j];
                scan_reg[(2*i)+1] = Addrb_r[j];
                end
              else if ((i >= 5) && (i < 8))
                begin
                j = i;
                scan_reg[2*i] = Addra_r[j];
                scan_reg[(2*i)+1] = Addrb_r[j];
                end
              else if ((i >= 8) && (i <= 9))
                begin
                j = i+2-1-9;
                scan_reg[2*i] = Addra_r[j];
                scan_reg[(2*i)+1] = Addrb_r[j];
                end
            end
	      
	    for (i = 0; i < BPW; i = i + 1)
	      begin
	        scan_reg[C1+2*i] = Wbtb_n_r[i];
	        scan_reg[C1+2*i+1] = Dinb_r[i];
	      end
	    for (i = 0; i < BPW; i = i + 1)
	      begin
	        douta[i] = scan_reg[C1+2*i+1];
	      end
	    sout = scan_reg[(2*BPW) + (2*SCAN_DEPTH_ADDR) + 1];
	end
     end
   endtask

   // Initialize entire memory to zero
   task initialize_memory;
      integer i;
      begin
       for (i = 0; i < WORDS; i = i + 1)
          begin
	   i_memArray[i] = 0;
          end
      end
   endtask

   task invalid_Csa_n_r;
      begin
         if (NO_WARNING == 0)
         if (scan_n === 1'b1 && clamp_mem === 1'b0 && slp_ret_n === 1'b1 && slp_nret_n === 1'b1)
         begin
           douta = {BPW{1'bx}};
         end
      end
   endtask

   // Invalidate scan registers 
   task invalidate_scan_registers;
      integer i;
      begin
	 for (i = 0; i < ((2*BPW) + (2*SCAN_DEPTH_ADDR) + 1) ; i = i + 1)
	   scan_reg[i] = 1'bx;
      end
   endtask

   task invalid_Csb_n_r;
      begin
         if (NO_WARNING == 0)
           $display(" %t : Warning on memory instance %m:: Write port chip select holding invalid value.", $time);
         if (scan_n === 1'b1 && clamp_mem === 1'b0 && slp_ret_n === 1'b1 && slp_nret_n === 1'b1)
          begin
	        if(^Addrb_rw === 1'bx)
		 invalidate_memory;
	        else
		 i_memArray[Addrb_rw] = {BPW{1'bx}};
           end
      end
   endtask

   task invalid_Addra_r;
      begin
         if (NO_WARNING == 0)
         $display(" %t : Warning on memory instance %m:: Read port address holding invalid value ", $time);
		douta = {BPW{1'bx}};
      end
   endtask

   task invalid_Addrb_r;
      begin
         if (NO_WARNING == 0)
         $display(" %t : Warning on memory instance %m:: Write port address holding invalid value", $time);
         invalidate_memory;
      end
   endtask

   task read;
      begin
         if(^Addra_rw === 1'bx)
           invalid_Addra_r;
         else if(^Addra_rw >= WORDS)
            begin
               if (NO_WARNING == 0)
                  $display(" %t : Warning on memory instance %m:: Address %d out of range ", $time, Addra_rw);
               douta = {BPW{1'bx}};
            end
         else
           douta = i_memArray[Addra_rw] ; 
        if (MEMORY_TRACE_LOG != "off")
          begin
             $fdisplay(log_file, " %0t (read) acc=%b addra=%b addrb=%b clamp_mem=%b clk=%b csa_n=%b csb_n=%b dinb=%b douta=%b scan_n=%b shift_n=%b sin=%b slp_nret_n=%b slp_ret_n=%b sout=%b %m", $time, acc, addra, addrb, clamp_mem, clk, csa_n, csb_n, dinb, douta, scan_n, shift_n, sin, slp_nret_n, slp_ret_n, sout);
             $fflush(log_file);
          end
      end
   endtask

   // Write into port B
   task write;
      begin
        if (MEMORY_TRACE_LOG != "off")
          begin
             $fdisplay(log_file, " %0t (write) acc=%b addra=%b addrb=%b clamp_mem=%b clk=%b csa_n=%b csb_n=%b dinb=%b douta=%b scan_n=%b shift_n=%b sin=%b slp_nret_n=%b slp_ret_n=%b sout=%b %m", $time, acc, addra, addrb, clamp_mem, clk, csa_n, csb_n, dinb, douta, scan_n, shift_n, sin, slp_nret_n, slp_ret_n, sout);
             $fflush(log_file);
          end
         if (^Addrb_rw === 1'bx)
             invalid_Addrb_r;
          else if(^Addrb_rw >= WORDS)
             begin
               if (NO_WARNING == 0)
                 $display(" %t : Warning on memory instance %m:: Address %d out of range ", $time, Addrb_rw);
             end
          else
            begin
              i_memArray[Addrb_rw] = Dinb_r;
            end
      end
   endtask

   task failure_inject_write;
     begin
       if (FAILURE_INJECT == 0)
	 begin
	 temp_write_failure_reg = temp_write_reg;
	 end
       else
	 begin
	  if(failed_io > BPW-1)
	   $display(" %t : Warning on memory instance %m :: failed_io %d is out of range", $time, failed_io);
	  else
	  begin
	   temp_write_failure_reg = temp_write_reg;
	   if(Addrb_rw == failed_addr)
	     begin
	      if (NO_WARNING == 0)
		begin
		$display(" %t : Warning on memory instance %m :: Failure Injection is ON and failed io is %b and failed addr is %h", $time, failed_io, failed_addr);
		end
	      temp_write_failure_reg[failed_io] = ~(temp_write_failure_reg[failed_io]);
	     end
	  end
	 end
     end
   endtask

   /**** Task definitions for use with VERA ****/
   task mem_write;
      input [ADDR_WIDTH - 1:0] address;
      input [BPW - 1:0] data;
      begin
	 if (address >= WORDS)
           begin
           if (NO_WARNING == 0)
	   $display(" %t : Warning on memory instance %m:: Address out of range ", $time);
           end
	 else if (^address === 1'bx)
	   begin
              if (NO_WARNING == 0)
	      $display(" %t : Error on memory instance %m:: Invalid address supplied to mem_write ", $time);
	   end
	 else
	   i_memArray[address] = data;
      end
   endtask

   task mem_read;
      input [ADDR_WIDTH - 1:0] address;
      output [BPW - 1:0] data;
      begin
	 if (address >= WORDS)
	   begin
              if (NO_WARNING == 0)
	      $display(" %t : Warning on memory instance %m:: Address out of range ", $time);
	      data = {BPW{1'bx}};
	   end
	 else if (^address === 1'bx)
	   begin
              if (NO_WARNING == 0)
	      $display(" %t : Error on memory instance %m:: Invalid address supplied to mem_read ", $time);
	      data = {BPW{1'bx}};
	   end
	 else
	   data = i_memArray[address];
      end
   endtask

   task mem_load;
      input [128 * 8 - 1:0] filename;
      begin
	 image_file = $fopen (filename, "r");
	 if (image_file == 0)
	   begin
	      $display(" %t : Error on memory instance %m:: Image file %0s cannot be opened. \n", $time, image_file);
	   end
	 $fclose (image_file);
	 $readmemh(filename, i_memArray);
      end
   endtask

   /***** Initial Block *****/
   initial
     begin
        $timeformat(-9, 0, " ns", 20);
        wait_period = 0;
        slp_min_period = 0;
        diff_time = 0;
        count = 0;
        current_time = 0;
        prev_time = 0;
        flag_tpd1 = 0;
        flag_tpd4 = 0;
        dummy_clock_reg = 0;
        #0 prev_slp_nret_n = slp_nret_n;
        $display("Memory instance %m created using QCmemmodel version 1.58 ");
        failed_io = FAILED_IO;
        failed_addr = FAILED_ADDR;
        // Check to see if trace log has been enabled for this instance
        // `ifndef _ESP_
        //$init_trace_1_58(NO_WARNING,NO_CORRUPT,IMAGE_FILE,MEMORY_TRACE_LOG);
        // `endif
        // See if a generic has been passed for image file loading
        case (filename)
           "NONE":
             begin
               $display("No image file associated with memory instance %m \n");

             end
           "ALL_ZERO":
             initialize_memory;
           "DEFAULT":
             begin
                // `ifndef _ESP_
                //$read_image_1_58;
                // `endif
                // If found, IMAGE_FILE is overwritten by path to image file
                if (IMAGE_FILE != "NULL")
                  begin
                     $display("Loading image file %0s for instance %m......", IMAGE_FILE);
                     $readmemh(IMAGE_FILE, i_memArray);
                     $display("done\n");
                  end
             end
           default:
             begin
              $display("Loading image file %0s for instance %m......", filename);
              $readmemh(filename, i_memArray);
             end
         endcase

         // If enabled, MEMORY_TRACE_LOG overwritten by name of trace log file
         if (MEMORY_TRACE_LOG == "off")
           $display ("No trace log associated with memory instance %m \n To enable trace log \'setenv MEMORY_TRACE_LOG on\'\n");
         else
           begin
              $display ("Enabling trace log for memory instance %m \n");
              log_file = $fopen(MEMORY_TRACE_LOG, "a");
              if (log_file == 0)
                begin
                   $display($time, " Error on memory instance %m:: File %s cannot be opened. \n", MEMORY_TRACE_LOG);
                end
              else
              // Trace file header information is printed
                begin
                   $fdisplay (log_file, "%m param_begin");
                   $fdisplay (log_file, "memory_name=cat_ram2p_half");
                   $fdisplay (log_file, "data_width=%0d", BPW);
                   $fdisplay (log_file, "addr_width=%0d", ADDR_WIDTH);
                   $fdisplay (log_file, "word_size=%0d", WORDS);
                   $fdisplay (log_file, "mux_option=4");
                   $fdisplay (log_file, "rising_edge=1");
                   $fdisplay (log_file, "param_end");
                   $fdisplay (log_file, "");
                   $fflush(log_file);
                end
           end
      end

   always @(csa_n, csb_n, addra, addrb, dinb, shift_n, scan_n, sin, scan_reg)
     begin
       get_wbtb_for_word;
       input_source_select;
     end

   always @(clk)
     begin
       if (wait_period == 1) 
	  begin
	     if ($time != 0) begin
               if (NO_WARNING == 0)
                 begin
	           $display (" %t : Error on memory instance %m:: Sleep violation, clk should be low for minimum 20ns after sleep de-assertion", $time);
                 end
	       invalidate_memory;// No need to invalidate scan registes since, in sleep mode scan registers are already invalidated 
             end
               douta = {BPW{1'bx}};
               sout = 1'bx;
	  end
	if (slp_min_period == 1) 
	  begin
	     if ($time != 0) begin
               if (NO_WARNING == 0)
                 begin
	           $display (" %t : Error on memory instance %m:: Sleep violation, clock should be zero for minimum 20ns after entering sleep mode", $time);
                 end
	       invalidate_memory;
             end
	       douta = {BPW{1'bx}};
	       sout = 1'bx;
	  end
	end

   always @(acc)
    $display(" %t : acc value has changed :: Value of acc %b in memory:%m", $time, acc);
   always @(acc, wait_period, slp_ret_n, slp_nret_n, clamp_mem)
     begin
      if ((wait_period == 0) &&((slp_ret_n === 1'b1) &&(slp_nret_n === 1'b1) && (clamp_mem === 1'b0)))
       begin
     if (^acc === 1'bx) begin
       valid_acc = 0;
       if ($time != 0) begin
         if (NO_WARNING == 0)
         begin
           $display(" %t : ERROR on memory instance %m :: Acc is x ", $time);
         end
         invalidate_memory;
       end
     end
     else begin
       valid_acc = 1;
     end
     end

      else begin
        valid_acc = 1;
      end
     end

   always @(posedge clk)
   begin
   count = count+1;

   if (count > 1 && slp_nret_n !== 1'b0 && slp_ret_n !== 1'b0 && clamp_mem === 1'b0) begin
     current_time = $time;
     diff_time = current_time - prev_time;
     if ((0 >= 20) || (diff_time >= 20)) begin
     diff_time = 20;
     end
     if ((0 > 0) && (0 < 20)) begin
     diff_time = 0 ;
     end
     prev_time = current_time;
    end
    else 
    begin
     current_time = $time;
     prev_time = current_time;
    end
   end

   always @(negedge clk)
     begin
       if(clamp_mem === 1'b0)
	     begin
	      if ((slp_ret_n === 1'b0) || (slp_nret_n === 1'b0))
	      begin
	      flag_tpd4 = 1;
	      flag_tpd4 = #5 0;
	      end
	      if ((slp_ret_n === 1'b1) && (slp_nret_n === 1'b1))
	      begin
	      flag_tpd1 = 1;
	      flag_tpd1 = #diff_time 0;
	      end
	     end
	    end

   always @(clk)
     begin
       casez ({prev_clk, clk})
         2'b00: ;
         2'b01:  begin 
           casez ({scan_n, shift_n})
             2'b0? ,
             2'b11: begin 
               register_inputs;
               register_rw_addr;
  // Adding constraint for cs_n to be high during dummy cycle after sleep
    		if (dummy_clock_reg === 1'b0 && slp_ret_n === 1'b1 && slp_nret_n === 1'b1 && clamp_mem === 1'b0 && scan_n === 1'b1 && wait_period === 1'b0)
    		begin
      		casez (Csb_n)
    	  		1'b0: begin
    	      		if (NO_WARNING == 0)
    	      		begin
    	      		$display("%t : Error on memory instance %m:: Chip select should be high for the 1st clock cycle (at posedge) after wakeup from sleep  !! ", $time);
    	      		end
    	   		if (NO_CORRUPT == 0)
    	   		begin
    	      		i_memArray[Addrb_r] = {BPW{1'bx}};
    	   		end
    	   		end
    	  		1'b1: ;
    	  		1'bx: ;
    	  		default: ;
      		endcase
      		casez (Csa_n)
    	  		1'b0: begin
    	      		if (NO_WARNING == 0)
    	      		begin
    	      		$display("%t : Warning on memory instance %m:: Chip select should be high for the 1st clock cycle (at posedge) after wakeup from sleep  !! ", $time);
    	      		end
    	      		douta = {BPW{1'bx}};
    	   		end
    	  		1'b1: ;
    	  		1'bx: ;
    	  		default: ;
      		endcase
    		end
               check_mode;
               mem_func;
               update_scan_reg;
             end 
             default: begin // This is illegal mode... 
		 casez ({clamp_mem, slp_ret_n, slp_nret_n}) // Here Giving Higher order of preference to clamp_mem and sleep than the Illegal mode.. 
		   3'b011:begin
                     invalidate_memory ;
                     invalidate_scan_registers ;
		     douta = {BPW{1'bx}}; 
		     sout = 1'bx;
                 end 
                 default: ;
               endcase
             end 
           endcase
	       // This is done after the update_scan_reg etc, hence for first clock cycle dummy_clock_reg will be 0 for wakeup. 
           if (wait_period == 0)
             begin
             if ((slp_ret_n === 1'b1) &&(slp_nret_n === 1'b1) && (clamp_mem === 1'b0))
               dummy_clock_reg  = 1;
             else
               dummy_clock_reg  = 0;
             end
	    end
         2'b10: ;
         2'b1x: ;
         default: ;
       endcase
       prev_clk = clk ;
     end

   always @(slp_ret_n, slp_nret_n, wait_period)
     begin
       casez ({clamp_mem, slp_ret_n, slp_nret_n, wait_period})
         4'b0x??: begin 
            if (NO_WARNING == 0)
              begin
                $display("  %t : Error on memory instance %m:: slp_ret_n holding invalid value ", $time);
              end
              if (slp_nret_n === 1'b0 )
	       begin
	        invalidate_memory_always;
	        douta = {BPW{1'b0}};
		sout = 1'b0;
  	       end
               if (slp_nret_n === 1'b1 || slp_nret_n === 1'bx)
	        begin
                 if (slp_nret_n === 1'bx)
                  begin
	           invalidate_memory;
                   if (NO_WARNING == 0)
                    begin
                    $display("  %t : Error on memory instance %m:: slp_ret_n holding invalid value ", $time);
                    end
                  end
	         douta = {BPW{1'bx}};
		 sout = 1'bx;
  	        end
	       invalidate_scan_registers;
               dummy_clock_reg = 0;
     	     end
         4'b0?x?: begin 
            if (NO_WARNING == 0)
              begin
                $display("  %t : Error on memory instance %m:: slp_nret_n holding invalid value ", $time);
              end
	        invalidate_memory;
	        invalidate_scan_registers;
                if (slp_ret_n === 1'b0 )
		 begin
		  douta = {BPW{1'b0}};
		  sout = 1'b0;
  		 end
                if (slp_ret_n === 1'b1 ||  slp_ret_n === 1'bx)
		 begin
                  if (NO_WARNING == 0 && slp_ret_n === 1'bx)
                    begin
                    $display("  %t : Warning on memory instance %m:: slp_ret_n holding invalid value ", $time);
                    end
		  douta = {BPW{1'bx}};
		  sout = 1'bx;
  		 end
            	dummy_clock_reg = 0;
     		end
         4'b00??: begin 
	          invalidate_scan_registers;
            	if (slp_nret_n === 1'b0 )
	          invalidate_memory_always;
                  if (slp_nret_n === 1'b1 || slp_nret_n === 1'bx)
		   begin
                    if (slp_nret_n === 1'bx)
                     begin
	              invalidate_memory;
                      if (NO_WARNING == 0)
                       begin
                       $display("  %t : Error on memory instance %m:: slp_ret_n holding invalid value ", $time);
                       end
                     end
                    end
            	douta = {BPW{1'b0}};
		sout = 1'b0;
            	dummy_clock_reg = 0;
     		end
         4'b0?0?: begin 
	    	  invalidate_memory_always;
	          invalidate_scan_registers;
            	  douta = {BPW{1'b0}};
		  sout = 1'b0;
            	  dummy_clock_reg = 0;
            	end
         4'b1???: begin 
	          invalidate_scan_registers;
            	douta = {BPW{1'b0}};
		sout = 1'b0;
            	dummy_clock_reg = 0;
     		end
         default: ;
       endcase
     end


   always @(negedge slp_ret_n, negedge slp_nret_n)
     begin
     if(clamp_mem === 1'b0)
     begin

     if (flag_tpd1 != 1'b0)
	begin
	 if (NO_WARNING == 0)
               begin
	         $display (" %t : Error on memory instance %m:: Sleep violation, clock should be zero for one clock cycle before sleep assertion", $time);
               end
	     invalidate_memory;
             douta = {BPW{1'bx}};
             sout = 1'bx;
	    end

     slp_min_period = 1;
     if ( clk !== 0 ) 
	  begin
	     if ($time != 0) begin
               if (NO_WARNING == 0)
                 begin
	           $display (" %t : Error on memory instance %m:: Sleep violation, clock should be low while sleep assertion ", $time);
                 end
	       invalidate_memory;
             end
               douta = {BPW{1'bx}};
               sout = 1'bx;
	    end
     slp_min_period = #20 0;
     end
     end


   always @(posedge slp_ret_n, posedge slp_nret_n)
     begin
      if(clamp_mem === 1'b0)
       begin
        if (slp_min_period == 1'b1)
	 begin
	  if (NO_WARNING == 0)
               begin
	         $display (" %t : Error on memory instance %m:: Sleep violation, minimum period of Sleep mode is 20ns", $time);
               end
	     invalidate_memory;
             douta = {BPW{1'bx}};
             sout = 1'bx;
	 end
    if (flag_tpd4 == 1'b1)
	 begin
	  if (NO_WARNING == 0)
               begin
	         $display (" %t : Error on memory instance %m:: Sleep violation, clock should be low for minimum 5ns before wake up", $time);
               end
	     invalidate_memory;
             douta = {BPW{1'bx}};
	     sout = 1'bx;
	 flag_tpd4 = 0; 
	 end
	if((slp_ret_n === 1'b1) && (slp_nret_n === 1'b1))
         begin
         douta = {BPW{1'bx}};
	 sout = 1'bx;
         end
	wait_period = 1;
	 if ( clk !== 0 ) 
	  begin
	     if ($time != 0) begin
               if (NO_WARNING == 0)
                 begin
	           $display (" %t :  Error on memory instance %m:: Sleep violation, clock should be low while sleep de-assertion", $time);
                 end
	       invalidate_memory;
	     end
               douta = {BPW{1'bx}};
	       sout = 1'bx;
	     end
	count = 0;
	wait_period = #20 0;
      end
     end


   always @(clamp_mem)
     begin
       casez ({prev_clamp_mem, clamp_mem})
         2'b00: ;
         2'b01: begin
	    clamp_violation_check;
	    prev_slp_nret_n = slp_nret_n;
	    douta = {BPW{1'b0}};
	    sout = 1'b0;
	    invalidate_scan_registers;
	    if(prev_slp_nret_n === 1'b0)
	    	begin
	        invalidate_memory_always;
	    	end
	    dummy_clock_reg = 0;
         end
         2'b10: begin
	    clamp_violation_check;
	    douta = {BPW{1'bx}};
	    sout = 1'bx;
	    if(slp_nret_n !== prev_slp_nret_n)
	    	begin
	    	 if (^prev_slp_nret_n !== 1'bx) begin
	    	   if(NO_WARNING == 0)
	    	   begin
	    	    $display (" %t : Error on memory instance %m:: Power Collapse violation, slp_nret_n changed during power collapse mode", $time);
	    	   end
	    	 invalidate_memory;
	    	 end
	    	end
         end
         2'b?x: begin
                    if (NO_WARNING == 0)
                     begin
                     $display("  %t : Warning on memory instance %m:: clamp_mem holding invalid value ", $time);
                     end
	    invalidate_memory;
	    invalidate_scan_registers;
	    douta = {BPW{1'bx}};
	    sout = 1'bx;
	    dummy_clock_reg = 0;
         end
         default: ;
       endcase
       prev_clamp_mem = clamp_mem;
     end

endmodule

`endif

 
`ifdef __cat_ram2p_half__ 

`else 

`define __cat_ram2p_half__ 

module cat_ram2p_half (
				acc,
				addra,
				addrb,
				clamp_mem,
				clk,
				csa_n,
				csb_n,
				dinb,
				douta,
				scan_n,
				shift_n,
				sin,
				slp_nret_n,
				slp_ret_n,
				sout
			);

  parameter filename = "DEFAULT" ;
  //parameter filename_size = 256 ;
  //parameter 0  = 0 ;
  parameter MEMORY_ACC_WIDTH  = 4;
  input [MEMORY_ACC_WIDTH-1:0] acc ;
  input [7:0] addra ;
  input [7:0] addrb ;
  input clamp_mem ;
  input clk ;
  input csa_n ;
  input csb_n ;
  input [63:0] dinb ;
  output [63:0] douta ;
  input scan_n ;
  input shift_n ;
  input sin ;
  input slp_nret_n ;
  input slp_ret_n ;
  output sout ;


  wire [3:0] i_acc ;
  wire [7:0] i_addra ;
  wire [7:0] i_addrb ;
  wire i_clamp_mem ;
  wire i_clk ;
  wire i_csa_n ;
  wire i_csb_n ;
  wire [63:0] i_dinb ;
  wire [63:0] i_douta ;
  wire i_scan_n ;
  wire i_shift_n ;
  wire i_sin ;
  wire i_slp_nret_n ;
  wire i_slp_ret_n ;
  wire i_sout ;


  assign douta = i_douta;
  assign sout = i_sout;


  buf #0 inst_acc [3:0] ( i_acc , acc ) ;
  buf #0 inst_addra [7:0] ( i_addra , addra ) ;
  buf #0 inst_addrb [7:0] ( i_addrb , addrb ) ;
  buf ( i_clamp_mem , clamp_mem ) ;
  buf ( i_clk , clk ) ;
  buf #0 ( i_csa_n , csa_n ) ;
  buf #0 ( i_csb_n , csb_n ) ;
  buf #0 inst_dinb [63:0] ( i_dinb , dinb ) ;
  buf #0 ( i_scan_n , scan_n ) ;
  buf #0 ( i_shift_n , shift_n ) ;
  buf #0 ( i_sin , sin ) ;
  buf ( i_slp_nret_n , slp_nret_n ) ;
  buf ( i_slp_ret_n , slp_ret_n ) ;

    core #(filename, 256) M1( 
    //core #(filename, filename_size) M1(
			.acc(i_acc),
			.addra(i_addra),
			.addrb(i_addrb),
			.clamp_mem(i_clamp_mem),
			.clk(i_clk),
			.csa_n(i_csa_n),
			.csb_n(i_csb_n),
			.dinb(i_dinb),
			.douta(i_douta),
			.scan_n(i_scan_n),
			.shift_n(i_shift_n),
			.sin(i_sin),
			.slp_nret_n(i_slp_nret_n),
			.slp_ret_n(i_slp_ret_n),
			.sout(i_sout)
			);

buf (delay_functional_mode ,scan_n );
and (scan_capture_mode ,!scan_n ,shift_n );
buf (scan_mode ,!scan_n );
and (scan_shift_mode ,!scan_n ,!shift_n );


specify
if (delay_functional_mode == 1'b1 )
( posedge clk *> ( douta +: M1.douta ) ) = ( 0 , 0 ) ;
if (scan_mode == 1'b1 )
( posedge clk *> ( douta +: M1.douta ) ) = ( 0 , 0 ) ;
if (scan_mode == 1'b1 )
( posedge clk *> ( sout +: M1.sout ) ) = ( 0 , 0 ) ;
$width ( posedge addra , 0 ) ;
$width ( negedge addra , 0 ) ;
$width ( posedge addrb , 0 ) ;
$width ( negedge addrb , 0 ) ;
$width ( posedge clk &&& (delay_functional_mode == 1'b1), 0 );
$width ( negedge clk &&& (delay_functional_mode == 1'b1), 0 );
$width ( posedge clk &&& (scan_mode == 1'b1), 0 );
$width ( negedge clk &&& (scan_mode == 1'b1), 0 );
$width ( posedge csa_n , 0 ) ;
$width ( negedge csa_n , 0 ) ;
$width ( posedge csb_n , 0 ) ;
$width ( negedge csb_n , 0 ) ;
$width ( posedge dinb , 0 ) ;
$width ( negedge dinb , 0 ) ;
$width ( posedge shift_n , 0 ) ;
$width ( negedge shift_n , 0 ) ;
$width ( posedge sin , 0 ) ;
$width ( negedge sin , 0 ) ;
$period ( posedge clk &&& (delay_functional_mode == 1'b1) , 0 );
$period ( posedge clk &&& (scan_mode == 1'b1) , 0 );
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , posedge addra &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , negedge addra &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , posedge addra &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , negedge addra &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , posedge addrb &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , negedge addrb &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , posedge addrb &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , negedge addrb &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , posedge csa_n &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , negedge csa_n &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , posedge csa_n &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , negedge csa_n &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , posedge csb_n &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , negedge csb_n &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , posedge csb_n &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , negedge csb_n &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , posedge dinb &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , negedge dinb &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , posedge dinb &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , negedge dinb &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_mode == 1'b1) , posedge shift_n &&& ( scan_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_mode == 1'b1) , negedge shift_n &&& ( scan_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_shift_mode == 1'b1) , posedge sin &&& ( scan_shift_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_shift_mode == 1'b1) , negedge sin &&& ( scan_shift_mode == 1'b1 ), 0 , 0 ) ;
$setuphold ( posedge clamp_mem, posedge slp_nret_n , 0 , 0 ) ; 
$setuphold ( posedge clamp_mem, negedge slp_nret_n , 0 , 0 ) ; 
$setuphold ( negedge clamp_mem, posedge slp_nret_n , 0 , 0 ) ; 
$setuphold ( negedge clamp_mem, negedge slp_nret_n , 0 , 0 ) ; 
$setuphold ( posedge clamp_mem, posedge slp_ret_n , 0 , 0 ) ; 
$setuphold ( posedge clamp_mem, negedge slp_ret_n , 0 , 0 ) ; 
$setuphold ( negedge clamp_mem, posedge slp_ret_n , 0 , 0 ) ; 
$setuphold ( negedge clamp_mem, negedge slp_ret_n , 0 , 0 ) ; 
endspecify
endmodule 

`endif 


//------> /hd/cad/mentor/2016.9/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v4.v 
module mgc_shift_r_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SIGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSIGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> /hd/cad/mentor/2016.9/Mgc_home/pkgs/siflibs/designcompiler/28nm.128x64.verilog.v 
// CONFIDENTIAL AND PROPRIETARY DATA OF QUALCOMM, INC. All Rights Reserved.
// Filename    	:    ram_lib.v
// Date        	:    Wed Mar 28 11:09:09 2018
// MTI .so file for sun32 and linux32 machines	:    /pkg/qcsw/memoryMagic2/QCmemmodel_28nm/1.58/pli/bin/qcmemmodel_pli_1_58.so
// MTI .so file for amd64 machine 		:    /pkg/qcsw/memoryMagic2/QCmemmodel_28nm/1.58/pli/bin/amd64/qcmemmodel_pli_1_58.so
// MTI .so file for sun64 machine 		:    /pkg/qcsw/memoryMagic2/QCmemmodel_28nm/1.58/pli/bin/sun64/qcmemmodel_pli_1_58.so
// PLI tab file 				:    /pkg/qcsw/memoryMagic2/QCmemmodel_28nm/1.58/pli/bin/qcmemmodel_pli_1_58.tab
// To refer the QCmemmodel FAQ page		:    http://qwiki.qualcomm.com/qct-ipmemory/QCmemmodel
// To refer the QCmemmodel User Guide		:    http://agiledocument.qualcomm.com/AgileDocument/spring/authorize?itemno=80-V9063-1&rev=YU
// ***please contact mem.help for any questions***


 
`ifdef __core__ 

`else 

`define __core__ 

module core (
				acc,
				addra,
				addrb,
				clamp_mem,
				clk,
				csa_n,
				csb_n,
				dinb,
				douta,
				scan_n,
				shift_n,
				sin,
				slp_nret_n,
				slp_ret_n,
				sout
			);
   // Parameter declarations
   parameter filename = "NONE";
   parameter filename_size = 128;
   parameter SCAN_DEPTH_ADDR = 9;
   parameter WORDS = 128;
   parameter ADDR_WIDTH = 7;
   parameter BPW = 64;
   parameter WORDX = {BPW{1'bx}};
   parameter FAILED_IO = 0;
   parameter FAILED_ADDR = 0;
   parameter SLEEP_TPD1 = 0;
   parameter ACC_DEBUG = 0;

   // Output and Input ports
   input	[3:0]	acc ;
   input	[6:0]	addra ;
   input	[6:0]	addrb ;
   input		clamp_mem ;
   input		clk ;
   input		csa_n ;
   input		csb_n ;
   input	[63:0]	dinb ;
   output	[63:0]	douta ;
   input		scan_n ;
   input		shift_n ;
   input		sin ;
   input		slp_nret_n ;
   input		slp_ret_n ;
   output		sout ;

   // Internal registers and memory array definitions
   reg                                                            prev_clk;
   reg [BPW - 1:0]                                                douta;
   reg                                                            sout;
   reg [BPW - 1:0]                                                Dinb;
   reg                                                            Csa_n;
   reg                                                            Csb_n;
   reg [BPW - 1:0]                                                Wbtb_n;
   reg [SCAN_DEPTH_ADDR :0]				          Addra;
   reg [SCAN_DEPTH_ADDR :0]				          Addrb;
   reg [SCAN_DEPTH_ADDR :0]				          Addra_r;
   reg [SCAN_DEPTH_ADDR :0]				          Addrb_r;
   reg [SCAN_DEPTH_ADDR :0]				          Addra_rw;
   reg [SCAN_DEPTH_ADDR :0]				          Addrb_rw;
   reg [BPW - 1:0]                                                Dinb_r;
   reg                                                            Csa_n_r;
   reg                                                            Csb_n_r;
   reg [BPW - 1:0]                                                Wbtb_n_r;
   reg                                                            wait_period;
   reg  	            			                  slp_min_period;
   reg                                                            flag_tpd4;
   reg                                                            flag_tpd1;
   reg [BPW - 1:0]                                                temp_write_reg;
   reg [BPW - 1:0]                                                temp_read_reg;
   reg [BPW - 1:0]                                                i_memArray [WORDS - 1:0];

   reg [BPW - 1:0]                                                wbtb_n;
   reg [2*BPW + 2*SCAN_DEPTH_ADDR + 1 : 0 ]            	  	  scan_reg;

   reg                                                            functional_mode;
   reg                                                            read_op;
   reg                                                            write_op;

   reg                                                            scan_op;

   reg                                                            dummy_clock_reg;
   reg                                                            prev_slp_nret_n;

   reg                                                            prev_clamp_mem;

   reg [8*filename_size - 1:0]                                    MEMORY_TRACE_LOG = "off";
   reg [8*filename_size - 1:0]                                    IMAGE_FILE = "NULL";
   reg                                                            NO_WARNING = 0;
   reg                                                            NO_CORRUPT = 0;
   reg                           		                  valid_acc = 0 ;
   integer                                                        log_file, image_file,count;
   reg                           		                  FAILURE_INJECT = 0 ;
   reg [BPW - 1:0] 	     	 				  temp_write_failure_reg;       // used for failure injection
   reg [5: 0]                           		          failed_io;
   reg [ADDR_WIDTH -1 : 0]                          failed_addr;
   time                                                        	prev_time, current_time, diff_time, sleep_time; 
   // Getting the memory modes
   task check_mode;
      begin
    // Adding waitperiod here to make sure nothing happens in wait period.. (dummy_clock_reg added for the same reason..) 
        functional_mode = scan_n & shift_n & dummy_clock_reg & ~clamp_mem & valid_acc & slp_ret_n & slp_nret_n;
        read_op = scan_n & shift_n & dummy_clock_reg & ~clamp_mem & valid_acc & slp_ret_n & slp_nret_n & (~Csa_n_r);
        write_op = scan_n & shift_n & dummy_clock_reg & ~clamp_mem & valid_acc  & slp_ret_n & slp_nret_n & (~Csb_n_r);
        scan_op = ~scan_n & ~clamp_mem & valid_acc & slp_ret_n & slp_nret_n;
      end
   endtask

   // Write all 1's into wbt_n for word writable memory
   task get_wbtb_for_word;
      // Loop Counter
      integer 	i;
      begin
         for (i = 0; i < BPW; i = i + 1)
             wbtb_n[i] = 1'b0;
      end
   endtask

   task get_Addra_Addrb;
      integer i;
      integer c;
      parameter last_addr = 9;
      begin
      c = 0;
      for(i = 2; i < 5; i = i+1)
      begin
      if(i == 2)
         begin
         Addra[i] = shift_n ? addra[i] : sin ;
         Addrb[i] = shift_n ? addrb[i] : scan_reg[(2*c)] ;
         c= c+1;
         end
      else if((i > 2) && (i < ADDR_WIDTH)) 
         begin
         Addra[i] = shift_n ? addra[i] : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? addrb[i] : scan_reg[(2*c)] ;
         c= c+1;
         end
      else
         begin
         Addra[i] = shift_n ? 1'b0 : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? 1'b0 : scan_reg[(2*c)] ;
         c= c+1;
         end
      end

      for(i = 8; i <= 9; i = i+1)
      begin
      if(i < ADDR_WIDTH)
         begin
         Addra[i] = shift_n ? addra[i] : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? addrb[i] : scan_reg[(2*c)] ;
         c= c+1;
         end
      else
         begin
         Addra[i] = shift_n ? 1'b0 : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? 1'b0 : scan_reg[(2*c)] ;
         c= c+1;
         end
      end

      for(i = 5; i < 8; i = i+1)
      begin
      if(i < ADDR_WIDTH)
         begin
         Addra[i] = shift_n ? addra[i] : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? addrb[i] : scan_reg[(2*c)] ;
         c= c+1;
         end
      else
         begin
         Addra[i] = shift_n ? 1'b0 : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? 1'b0 : scan_reg[(2*c)] ;
         c= c+1;
         end
      end

      for(i = 0; i < 2; i = i+1)
      begin
      if(i < ADDR_WIDTH)
         begin
         Addra[i] = shift_n ? addra[i] : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? addrb[i] : scan_reg[(2*c)] ;
         c= c+1;
         end
      else
         begin
         Addra[i] = shift_n ? 1'b0 : scan_reg[(2*c)-1] ;
         Addrb[i] = shift_n ? 1'b0 : scan_reg[(2*c)] ;
         c= c+1;
         end
      end
   end
   endtask

   task get_Csa_n;
      begin
    Csa_n = csa_n ;
      end
   endtask

   task get_Csb_n;
      begin
    Csb_n = csb_n ;
      end
   endtask

   // Getting Din through scan logic
   // The selection is between previous scan register( width = addr_width + 1; ie 0 to addr_width; din[0] has to choose between  scan reg[addr_width] and normal din logic.  
   task get_Wbtn_n_Dinb;
      integer i;
      integer j;
      parameter C1 = 2 * SCAN_DEPTH_ADDR + 2;
      begin
	 for (i = 0; i < BPW; i = i + 1)
	   begin
	       Wbtb_n[i] = shift_n ? wbtb_n[i] : scan_reg[C1+(2*i) -1] ;
	       Dinb[i] = shift_n ? dinb[i] : scan_reg[C1+(2*i)] ;
	   end
      end
   endtask

   // Write into specified bits alone
   task bit_wise_write;
      integer i;
      begin
      for (i = 0; i < BPW; i = i + 1)
        if (!Wbtb_n_r[i])
 	 temp_write_reg[i] = Dinb_r[i];
      end
   endtask

   // Select between BIST and normal inputs
   task input_source_select;
      begin
      get_Addra_Addrb ;
      get_Csa_n ;
      get_Csb_n ;
      get_Wbtn_n_Dinb ;
      end
   endtask

   // Register inputs
   task register_inputs;
      begin
	Dinb_r     = Dinb ; 
	Addra_r    = Addra ; 
	Addrb_r    = Addrb ; 
        Wbtb_n_r   = Wbtb_n ; 
        Csa_n_r    = Csa_n ; 
        Csb_n_r    = Csb_n ; 
      end
   endtask

   // Register read/write address
   task register_rw_addr;
     parameter MSB1 = 9;
     parameter MSB2 = 8;
       begin
	 Addra_rw    = Addra_r ; 
	 Addrb_rw    = Addrb_r ; 
      end
   endtask

   // Invalidate entire memory
   task invalidate_memory;
      integer i;
      begin
         if (NO_CORRUPT == 0)
           begin
            if (NO_WARNING == 0)
              begin
              $display(" %t : Memory instance %m:: Invalidating memory contents ", $time);
              end
	    for (i = 0; i < WORDS; i = i + 1)
	       begin
	        i_memArray[i] = WORDX;
	       end
      end
         else
           begin
             if (NO_WARNING == 0)
               begin
                 $display("%t : Warning on memory instance %m:: NO_CORRUPT Flag is set and hence invalid inputs wont corrupt the memory !! ", $time);
               end
          end
      end
   endtask

   // Invalidate entire memory for sleep no retention
   task invalidate_memory_always;
      integer i;
      begin
	 if (NO_CORRUPT == 0)
	   begin
	    if (NO_WARNING == 0)
	      begin
	      $display(" %t : Memory instance %m:: Invalidating memory contents ", $time);
	      end
	    for (i = 0; i < WORDS; i = i + 1)
	       begin
	        i_memArray[i] = WORDX;
	       end
	   end
	 else
	   begin
	     if (NO_WARNING == 0)
	       begin
		 $display("%t : Warning on memory instance %m:: NO_CORRUPT Flag is set and hence sleep no retention mode wont corrupt the memory !! ", $time);
	       end
	   end
      end
   endtask

   // Clk and slp_ret_n should be zero when the clamp_mem is asserted or de-asserted
   task clamp_violation_check;
      begin
         if ((slp_ret_n !== 1'b0) && (slp_nret_n !== 1'b0))
           begin
             if (NO_WARNING == 0)
               begin
                 $display("%t : Error on memory instance %m:: Power Collapse Violation. slp_ret_n should be low ", $time);
               end
             invalidate_memory;
          end
      end
   endtask

   // memory functional cycle 
   task mem_func;
      begin
        if(wait_period == 0)
          begin
           if ( read_op == 1 )
              read ;
           if ( write_op == 1 )
              write ;
           if ((Csa_n_r === 1'bx) && ( functional_mode == 1 ))
              invalid_Csa_n_r ;
           if ((Csb_n_r === 1'bx) && ( functional_mode == 1 ))
              invalid_Csb_n_r ;
          end
      end
   endtask

   // Updating the scan chain
   task update_scan_reg;
     integer i ;
     integer j ;
     parameter C1 = 2*SCAN_DEPTH_ADDR + 2 ;
     begin
        if (scan_op == 1)
        begin
	    for (i = 0; i <= SCAN_DEPTH_ADDR; i = i + 1)
            begin
              if (i < 3)
                begin
                j = 2+i;
                scan_reg[2*i] = Addra_r[j];
                scan_reg[(2*i)+1] = Addrb_r[j];
                end
              else if ((i == 3) || (i == 4))
                begin
                j = 9-4+i;
                scan_reg[2*i] = Addra_r[j];
                scan_reg[(2*i)+1] = Addrb_r[j];
                end
              else if ((i >= 5) && (i < 8))
                begin
                j = i;
                scan_reg[2*i] = Addra_r[j];
                scan_reg[(2*i)+1] = Addrb_r[j];
                end
              else if ((i >= 8) && (i <= 9))
                begin
                j = i+2-1-9;
                scan_reg[2*i] = Addra_r[j];
                scan_reg[(2*i)+1] = Addrb_r[j];
                end
            end
	      
	    for (i = 0; i < BPW; i = i + 1)
	      begin
	        scan_reg[C1+2*i] = Wbtb_n_r[i];
	        scan_reg[C1+2*i+1] = Dinb_r[i];
	      end
	    for (i = 0; i < BPW; i = i + 1)
	      begin
	        douta[i] = scan_reg[C1+2*i+1];
	      end
	    sout = scan_reg[(2*BPW) + (2*SCAN_DEPTH_ADDR) + 1];
	end
     end
   endtask

   // Initialize entire memory to zero
   task initialize_memory;
      integer i;
      begin
       for (i = 0; i < WORDS; i = i + 1)
          begin
	   i_memArray[i] = 0;
          end
      end
   endtask

   task invalid_Csa_n_r;
      begin
         if (NO_WARNING == 0)
         if (scan_n === 1'b1 && clamp_mem === 1'b0 && slp_ret_n === 1'b1 && slp_nret_n === 1'b1)
         begin
           douta = WORDX;
         end
      end
   endtask

   // Invalidate scan registers 
   task invalidate_scan_registers;
      integer i;
      begin
	 for (i = 0; i < ((2*BPW) + (2*SCAN_DEPTH_ADDR) + 1) ; i = i + 1)
	   scan_reg[i] = 1'bx;
      end
   endtask

   task invalid_Csb_n_r;
      begin
         if (NO_WARNING == 0)
           $display(" %t : Warning on memory instance %m:: Write port chip select holding invalid value.", $time);
         if (scan_n === 1'b1 && clamp_mem === 1'b0 && slp_ret_n === 1'b1 && slp_nret_n === 1'b1)
          begin
	        if(^Addrb_rw === 1'bx)
		 invalidate_memory;
	        else
		 i_memArray[Addrb_rw] = WORDX;
           end
      end
   endtask

   task invalid_Addra_r;
      begin
         if (NO_WARNING == 0)
         $display(" %t : Warning on memory instance %m:: Read port address holding invalid value ", $time);
		douta = WORDX;
      end
   endtask

   task invalid_Addrb_r;
      begin
         if (NO_WARNING == 0)
         $display(" %t : Warning on memory instance %m:: Write port address holding invalid value", $time);
         invalidate_memory;
      end
   endtask

   task read;
      begin
         if(^Addra_rw === 1'bx)
           invalid_Addra_r;
         else if(^Addra_rw >= WORDS)
            begin
               if (NO_WARNING == 0)
                  $display(" %t : Warning on memory instance %m:: Address %d out of range ", $time, Addra_rw);
               douta = WORDX;
            end
         else
           douta = i_memArray[Addra_rw] ; 
        if (MEMORY_TRACE_LOG != "off")
          begin
             $fdisplay(log_file, " %0t (read) acc=%b addra=%b addrb=%b clamp_mem=%b clk=%b csa_n=%b csb_n=%b dinb=%b douta=%b scan_n=%b shift_n=%b sin=%b slp_nret_n=%b slp_ret_n=%b sout=%b %m", $time, acc, addra, addrb, clamp_mem, clk, csa_n, csb_n, dinb, douta, scan_n, shift_n, sin, slp_nret_n, slp_ret_n, sout);
             $fflush(log_file);
          end
      end
   endtask

   // Write into port B
   task write;
      begin
        if (MEMORY_TRACE_LOG != "off")
          begin
             $fdisplay(log_file, " %0t (write) acc=%b addra=%b addrb=%b clamp_mem=%b clk=%b csa_n=%b csb_n=%b dinb=%b douta=%b scan_n=%b shift_n=%b sin=%b slp_nret_n=%b slp_ret_n=%b sout=%b %m", $time, acc, addra, addrb, clamp_mem, clk, csa_n, csb_n, dinb, douta, scan_n, shift_n, sin, slp_nret_n, slp_ret_n, sout);
             $fflush(log_file);
          end
         if (^Addrb_rw === 1'bx)
             invalid_Addrb_r;
          else if(^Addrb_rw >= WORDS)
             begin
               if (NO_WARNING == 0)
                 $display(" %t : Warning on memory instance %m:: Address %d out of range ", $time, Addrb_rw);
             end
          else
            begin
              i_memArray[Addrb_rw] = Dinb_r;
            end
      end
   endtask

   task failure_inject_write;
     begin
       if (FAILURE_INJECT == 0)
	 begin
	 temp_write_failure_reg = temp_write_reg;
	 end
       else
	 begin
	  if(failed_io > BPW-1)
	   $display(" %t : Warning on memory instance %m :: failed_io %d is out of range", $time, failed_io);
	  else
	  begin
	   temp_write_failure_reg = temp_write_reg;
	   if(Addrb_rw == failed_addr)
	     begin
	      if (NO_WARNING == 0)
		begin
		$display(" %t : Warning on memory instance %m :: Failure Injection is ON and failed io is %b and failed addr is %h", $time, failed_io, failed_addr);
		end
	      temp_write_failure_reg[failed_io] = ~(temp_write_failure_reg[failed_io]);
	     end
	  end
	 end
     end
   endtask

   /**** Task definitions for use with VERA ****/
   task mem_write;
      input [ADDR_WIDTH - 1:0] address;
      input [BPW - 1:0] data;
      begin
	 if (address >= WORDS)
           begin
           if (NO_WARNING == 0)
	   $display(" %t : Warning on memory instance %m:: Address out of range ", $time);
           end
	 else if (^address === 1'bx)
	   begin
              if (NO_WARNING == 0)
	      $display(" %t : Error on memory instance %m:: Invalid address supplied to mem_write ", $time);
	   end
	 else
	   i_memArray[address] = data;
      end
   endtask

   task mem_read;
      input [ADDR_WIDTH - 1:0] address;
      output [BPW - 1:0] data;
      begin
	 if (address >= WORDS)
	   begin
              if (NO_WARNING == 0)
	      $display(" %t : Warning on memory instance %m:: Address out of range ", $time);
	      data = WORDX;
	   end
	 else if (^address === 1'bx)
	   begin
              if (NO_WARNING == 0)
	      $display(" %t : Error on memory instance %m:: Invalid address supplied to mem_read ", $time);
	      data = WORDX;
	   end
	 else
	   data = i_memArray[address];
      end
   endtask

   task mem_load;
      input [filename_size * 8 - 1:0] filename;
      begin
	 image_file = $fopen (filename, "r");
	 if (image_file == 0)
	   begin
	      $display(" %t : Error on memory instance %m:: Image file %0s cannot be opened. \n", $time, image_file);
	   end
	 $fclose (image_file);
	 $readmemh(filename, i_memArray);
      end
   endtask

   /***** Initial Block *****/
   initial
     begin
        $timeformat(-9, 0, " ns", 20);
        wait_period = 0;
        slp_min_period = 0;
        diff_time = 0;
        count = 0;
        current_time = 0;
        prev_time = 0;
        flag_tpd1 = 0;
        flag_tpd4 = 0;
        dummy_clock_reg = 0;
        #0 prev_slp_nret_n = slp_nret_n;
        $display("Memory instance %m created using QCmemmodel version 1.58 ");
        failed_io = FAILED_IO;
        failed_addr = FAILED_ADDR;
        // Check to see if trace log has been enabled for this instance
        // `ifndef _ESP_
        $init_trace_1_58(NO_WARNING,NO_CORRUPT,IMAGE_FILE,MEMORY_TRACE_LOG);
        // `endif
        // See if a generic has been passed for image file loading
        case (filename)
           "NONE":
             begin
               $display("No image file associated with memory instance %m \n");

             end
           "ALL_ZERO":
             initialize_memory;
           "DEFAULT":
             begin
                // `ifndef _ESP_
                $read_image_1_58;
                // `endif
                // If found, IMAGE_FILE is overwritten by path to image file
                if (IMAGE_FILE != "NULL")
                  begin
                     $display("Loading image file %0s for instance %m......", IMAGE_FILE);
                     $readmemh(IMAGE_FILE, i_memArray);
                     $display("done\n");
                  end
             end
           default:
             begin
              $display("Loading image file %0s for instance %m......", filename);
              $readmemh(filename, i_memArray);
             end
         endcase

         // If enabled, MEMORY_TRACE_LOG overwritten by name of trace log file
         if (MEMORY_TRACE_LOG == "off")
           $display ("No trace log associated with memory instance %m \n To enable trace log \'setenv MEMORY_TRACE_LOG on\'\n");
         else
           begin
              $display ("Enabling trace log for memory instance %m \n");
              log_file = $fopen(MEMORY_TRACE_LOG, "a");
              if (log_file == 0)
                begin
                   $display($time, " Error on memory instance %m:: File %s cannot be opened. \n", MEMORY_TRACE_LOG);
                end
              else
              // Trace file header information is printed
                begin
                   $fdisplay (log_file, "%m param_begin");
                   $fdisplay (log_file, "memory_name=cat_ram2p_half_128x64");
                   $fdisplay (log_file, "data_width=%0d", BPW);
                   $fdisplay (log_file, "addr_width=%0d", ADDR_WIDTH);
                   $fdisplay (log_file, "word_size=%0d", WORDS);
                   $fdisplay (log_file, "mux_option=4");
                   $fdisplay (log_file, "rising_edge=1");
                   $fdisplay (log_file, "param_end");
                   $fdisplay (log_file, "");
                   $fflush(log_file);
                end
           end
      end

   always @(csa_n, csb_n, addra, addrb, dinb, shift_n, scan_n, sin, scan_reg)
     begin
       get_wbtb_for_word;
       input_source_select;
     end

   always @(clk)
     begin
       if (wait_period == 1) 
	  begin
	     if ($time != 0) begin
               if (NO_WARNING == 0)
                 begin
	           $display (" %t : Error on memory instance %m:: Sleep violation, clk should be low for minimum 20ns after sleep de-assertion", $time);
                 end
	       invalidate_memory;// No need to invalidate scan registes since, in sleep mode scan registers are already invalidated 
             end
               douta = WORDX;
               sout = 1'bx;
	  end
	if (slp_min_period == 1) 
	  begin
	     if ($time != 0) begin
               if (NO_WARNING == 0)
                 begin
	           $display (" %t : Error on memory instance %m:: Sleep violation, clock should be zero for minimum 20ns after entering sleep mode", $time);
                 end
	       invalidate_memory;
             end
	       douta = WORDX;
	       sout = 1'bx;
	  end
	end

   always @(acc)
    $display(" %t : acc value has changed :: Value of acc %b in memory:%m", $time, acc);
   always @(acc, wait_period, slp_ret_n, slp_nret_n, clamp_mem)
     begin
      if ((wait_period == 0) &&((slp_ret_n === 1'b1) &&(slp_nret_n === 1'b1) && (clamp_mem === 1'b0)))
       begin
     if (^acc === 1'bx) begin
       valid_acc = 0;
       if ($time != 0) begin
         if (NO_WARNING == 0)
         begin
           $display(" %t : ERROR on memory instance %m :: Acc is x ", $time);
         end
         invalidate_memory;
       end
     end
     else begin
       valid_acc = 1;
     end
     end

      else begin
        valid_acc = 1;
      end
     end

   always @(posedge clk)
   begin
   count = count+1;

   if (count > 1 && slp_nret_n !== 1'b0 && slp_ret_n !== 1'b0 && clamp_mem === 1'b0) begin
     current_time = $time;
     diff_time = current_time - prev_time;
     if ((SLEEP_TPD1 >= 20) || (diff_time >= 20)) begin
     diff_time = 20;
     end
     if ((SLEEP_TPD1 > 0) && (SLEEP_TPD1 < 20)) begin
     diff_time = SLEEP_TPD1 ;
     end
     prev_time = current_time;
    end
    else 
    begin
     current_time = $time;
     prev_time = current_time;
    end
   end

   always @(negedge clk)
     begin
       if(clamp_mem === 1'b0)
	     begin
	      if ((slp_ret_n === 1'b0) || (slp_nret_n === 1'b0))
	      begin
	      flag_tpd4 = 1;
	      flag_tpd4 = #5 0;
	      end
	      if ((slp_ret_n === 1'b1) && (slp_nret_n === 1'b1))
	      begin
	      flag_tpd1 = 1;
	      flag_tpd1 = #diff_time 0;
	      end
	     end
	    end

   always @(clk)
     begin
       casez ({prev_clk, clk})
         2'b00: ;
         2'b01:  begin 
           casez ({scan_n, shift_n})
             2'b0? ,
             2'b11: begin 
               register_inputs;
               register_rw_addr;
  // Adding constraint for cs_n to be high during dummy cycle after sleep
    		if (dummy_clock_reg === 1'b0 && slp_ret_n === 1'b1 && slp_nret_n === 1'b1 && clamp_mem === 1'b0 && scan_n === 1'b1 && wait_period === 1'b0)
    		begin
      		casez (Csb_n)
    	  		1'b0: begin
    	      		if (NO_WARNING == 0)
    	      		begin
    	      		$display("%t : Error on memory instance %m:: Chip select should be high for the 1st clock cycle (at posedge) after wakeup from sleep  !! ", $time);
    	      		end
    	   		if (NO_CORRUPT == 0)
    	   		begin
    	      		i_memArray[Addrb_r] = WORDX;
    	   		end
    	   		end
    	  		1'b1: ;
    	  		1'bx: ;
    	  		default: ;
      		endcase
      		casez (Csa_n)
    	  		1'b0: begin
    	      		if (NO_WARNING == 0)
    	      		begin
    	      		$display("%t : Warning on memory instance %m:: Chip select should be high for the 1st clock cycle (at posedge) after wakeup from sleep  !! ", $time);
    	      		end
    	      		douta = WORDX;
    	   		end
    	  		1'b1: ;
    	  		1'bx: ;
    	  		default: ;
      		endcase
    		end
               check_mode;
               mem_func;
               update_scan_reg;
             end 
             default: begin // This is illegal mode... 
		 casez ({clamp_mem, slp_ret_n, slp_nret_n}) // Here Giving Higher order of preference to clamp_mem and sleep than the Illegal mode.. 
		   3'b011:begin
                     invalidate_memory ;
                     invalidate_scan_registers ;
		     douta = WORDX; 
		     sout = 1'bx;
                 end 
                 default: ;
               endcase
             end 
           endcase
	       // This is done after the update_scan_reg etc, hence for first clock cycle dummy_clock_reg will be 0 for wakeup. 
           if (wait_period == 0)
             begin
             if ((slp_ret_n === 1'b1) &&(slp_nret_n === 1'b1) && (clamp_mem === 1'b0))
               dummy_clock_reg  = 1;
             else
               dummy_clock_reg  = 0;
             end
	    end
         2'b10: ;
         2'b1x: ;
         default: ;
       endcase
       prev_clk = clk ;
     end

   always @(slp_ret_n, slp_nret_n, wait_period)
     begin
       casez ({clamp_mem, slp_ret_n, slp_nret_n, wait_period})
         4'b0x??: begin 
            if (NO_WARNING == 0)
              begin
                $display("  %t : Error on memory instance %m:: slp_ret_n holding invalid value ", $time);
              end
              if (slp_nret_n === 1'b0 )
	       begin
	        invalidate_memory_always;
	        douta = {BPW{1'b0}};
		sout = 1'b0;
  	       end
               if (slp_nret_n === 1'b1 || slp_nret_n === 1'bx)
	        begin
                 if (slp_nret_n === 1'bx)
                  begin
	           invalidate_memory;
                   if (NO_WARNING == 0)
                    begin
                    $display("  %t : Error on memory instance %m:: slp_ret_n holding invalid value ", $time);
                    end
                  end
	         douta = WORDX;
		 sout = 1'bx;
  	        end
	       invalidate_scan_registers;
               dummy_clock_reg = 0;
     	     end
         4'b0?x?: begin 
            if (NO_WARNING == 0)
              begin
                $display("  %t : Error on memory instance %m:: slp_nret_n holding invalid value ", $time);
              end
	        invalidate_memory;
	        invalidate_scan_registers;
                if (slp_ret_n === 1'b0 )
		 begin
		  douta = {BPW{1'b0}};
		  sout = 1'b0;
  		 end
                if (slp_ret_n === 1'b1 ||  slp_ret_n === 1'bx)
		 begin
                  if (NO_WARNING == 0 && slp_ret_n === 1'bx)
                    begin
                    $display("  %t : Warning on memory instance %m:: slp_ret_n holding invalid value ", $time);
                    end
		  douta = WORDX;
		  sout = 1'bx;
  		 end
            	dummy_clock_reg = 0;
     		end
         4'b00??: begin 
	          invalidate_scan_registers;
            	if (slp_nret_n === 1'b0 )
	          invalidate_memory_always;
                  if (slp_nret_n === 1'b1 || slp_nret_n === 1'bx)
		   begin
                    if (slp_nret_n === 1'bx)
                     begin
	              invalidate_memory;
                      if (NO_WARNING == 0)
                       begin
                       $display("  %t : Error on memory instance %m:: slp_ret_n holding invalid value ", $time);
                       end
                     end
                    end
            	douta = {BPW{1'b0}};
		sout = 1'b0;
            	dummy_clock_reg = 0;
     		end
         4'b0?0?: begin 
	    	  invalidate_memory_always;
	          invalidate_scan_registers;
            	  douta = {BPW{1'b0}};
		  sout = 1'b0;
            	  dummy_clock_reg = 0;
            	end
         4'b1???: begin 
	          invalidate_scan_registers;
            	douta = {BPW{1'b0}};
		sout = 1'b0;
            	dummy_clock_reg = 0;
     		end
         default: ;
       endcase
     end


   always @(negedge slp_ret_n, negedge slp_nret_n)
     begin
     if(clamp_mem === 1'b0)
     begin

     if (flag_tpd1 != 1'b0)
	begin
	 if (NO_WARNING == 0)
               begin
	         $display (" %t : Error on memory instance %m:: Sleep violation, clock should be zero for one clock cycle before sleep assertion", $time);
               end
	     invalidate_memory;
             douta = WORDX;
             sout = 1'bx;
	    end

     slp_min_period = 1;
     if ( clk !== 0 ) 
	  begin
	     if ($time != 0) begin
               if (NO_WARNING == 0)
                 begin
	           $display (" %t : Error on memory instance %m:: Sleep violation, clock should be low while sleep assertion ", $time);
                 end
	       invalidate_memory;
             end
               douta = WORDX;
               sout = 1'bx;
	    end
     slp_min_period = #20 0;
     end
     end


   always @(posedge slp_ret_n, posedge slp_nret_n)
     begin
      if(clamp_mem === 1'b0)
       begin
        if (slp_min_period == 1'b1)
	 begin
	  if (NO_WARNING == 0)
               begin
	         $display (" %t : Error on memory instance %m:: Sleep violation, minimum period of Sleep mode is 20ns", $time);
               end
	     invalidate_memory;
             douta = WORDX;
             sout = 1'bx;
	 end
    if (flag_tpd4 == 1'b1)
	 begin
	  if (NO_WARNING == 0)
               begin
	         $display (" %t : Error on memory instance %m:: Sleep violation, clock should be low for minimum 5ns before wake up", $time);
               end
	     invalidate_memory;
             douta = WORDX;
	     sout = 1'bx;
	 flag_tpd4 = 0; 
	 end
	if((slp_ret_n === 1'b1) && (slp_nret_n === 1'b1))
         begin
         douta = WORDX;
	 sout = 1'bx;
         end
	wait_period = 1;
	 if ( clk !== 0 ) 
	  begin
	     if ($time != 0) begin
               if (NO_WARNING == 0)
                 begin
	           $display (" %t :  Error on memory instance %m:: Sleep violation, clock should be low while sleep de-assertion", $time);
                 end
	       invalidate_memory;
	     end
               douta = WORDX;
	       sout = 1'bx;
	     end
	count = 0;
	wait_period = #20 0;
      end
     end


   always @(clamp_mem)
     begin
       casez ({prev_clamp_mem, clamp_mem})
         2'b00: ;
         2'b01: begin
	    clamp_violation_check;
	    prev_slp_nret_n = slp_nret_n;
	    douta = {BPW{1'b0}};
	    sout = 1'b0;
	    invalidate_scan_registers;
	    if(prev_slp_nret_n === 1'b0)
	    	begin
	        invalidate_memory_always;
	    	end
	    dummy_clock_reg = 0;
         end
         2'b10: begin
	    clamp_violation_check;
	    douta = WORDX;
	    sout = 1'bx;
	    if(slp_nret_n !== prev_slp_nret_n)
	    	begin
	    	 if (^prev_slp_nret_n !== 1'bx) begin
	    	   if(NO_WARNING == 0)
	    	   begin
	    	    $display (" %t : Error on memory instance %m:: Power Collapse violation, slp_nret_n changed during power collapse mode", $time);
	    	   end
	    	 invalidate_memory;
	    	 end
	    	end
         end
         2'b?x: begin
                    if (NO_WARNING == 0)
                     begin
                     $display("  %t : Warning on memory instance %m:: clamp_mem holding invalid value ", $time);
                     end
	    invalidate_memory;
	    invalidate_scan_registers;
	    douta = WORDX;
	    sout = 1'bx;
	    dummy_clock_reg = 0;
         end
         default: ;
       endcase
       prev_clamp_mem = clamp_mem;
     end

endmodule

`endif

 
`ifdef __cat_ram2p_half_128x64__ 

`else 

`define __cat_ram2p_half_128x64__ 

module cat_ram2p_half_128x64 (
				acc,
				addra,
				addrb,
				clamp_mem,
				clk,
				csa_n,
				csb_n,
				dinb,
				douta,
				scan_n,
				shift_n,
				sin,
				slp_nret_n,
				slp_ret_n,
				sout
			);

  parameter filename = "DEFAULT" ;
  parameter filename_size = 256 ;
  parameter VLOG_DELAY  = 0 ;
  parameter MEMORY_ACC_WIDTH  = 4;
  input [MEMORY_ACC_WIDTH-1:0] acc ;
  input [6:0] addra ;
  input [6:0] addrb ;
  input clamp_mem ;
  input clk ;
  input csa_n ;
  input csb_n ;
  input [63:0] dinb ;
  output [63:0] douta ;
  input scan_n ;
  input shift_n ;
  input sin ;
  input slp_nret_n ;
  input slp_ret_n ;
  output sout ;


  wire [3:0] i_acc ;
  wire [6:0] i_addra ;
  wire [6:0] i_addrb ;
  wire i_clamp_mem ;
  wire i_clk ;
  wire i_csa_n ;
  wire i_csb_n ;
  wire [63:0] i_dinb ;
  wire [63:0] i_douta ;
  wire i_scan_n ;
  wire i_shift_n ;
  wire i_sin ;
  wire i_slp_nret_n ;
  wire i_slp_ret_n ;
  wire i_sout ;


  assign douta = i_douta;
  assign sout = i_sout;


  buf #VLOG_DELAY inst_acc [3:0] ( i_acc , acc ) ;
  buf #VLOG_DELAY inst_addra [6:0] ( i_addra , addra ) ;
  buf #VLOG_DELAY inst_addrb [6:0] ( i_addrb , addrb ) ;
  buf ( i_clamp_mem , clamp_mem ) ;
  buf ( i_clk , clk ) ;
  buf #VLOG_DELAY ( i_csa_n , csa_n ) ;
  buf #VLOG_DELAY ( i_csb_n , csb_n ) ;
  buf #VLOG_DELAY inst_dinb [63:0] ( i_dinb , dinb ) ;
  buf #VLOG_DELAY ( i_scan_n , scan_n ) ;
  buf #VLOG_DELAY ( i_shift_n , shift_n ) ;
  buf #VLOG_DELAY ( i_sin , sin ) ;
  buf ( i_slp_nret_n , slp_nret_n ) ;
  buf ( i_slp_ret_n , slp_ret_n ) ;


    core #(filename, filename_size) M1(
			.acc(i_acc),
			.addra(i_addra),
			.addrb(i_addrb),
			.clamp_mem(i_clamp_mem),
			.clk(i_clk),
			.csa_n(i_csa_n),
			.csb_n(i_csb_n),
			.dinb(i_dinb),
			.douta(i_douta),
			.scan_n(i_scan_n),
			.shift_n(i_shift_n),
			.sin(i_sin),
			.slp_nret_n(i_slp_nret_n),
			.slp_ret_n(i_slp_ret_n),
			.sout(i_sout)
			);

buf (delay_functional_mode ,scan_n );
and (scan_capture_mode ,!scan_n ,shift_n );
buf (scan_mode ,!scan_n );
and (scan_shift_mode ,!scan_n ,!shift_n );


specify
if (delay_functional_mode == 1'b1 )
( posedge clk *> ( douta +: M1.douta ) ) = ( 0 , 0 ) ;
if (scan_mode == 1'b1 )
( posedge clk *> ( douta +: M1.douta ) ) = ( 0 , 0 ) ;
if (scan_mode == 1'b1 )
( posedge clk *> ( sout +: M1.sout ) ) = ( 0 , 0 ) ;
$width ( posedge addra , 0 ) ;
$width ( negedge addra , 0 ) ;
$width ( posedge addrb , 0 ) ;
$width ( negedge addrb , 0 ) ;
$width ( posedge clk &&& (delay_functional_mode == 1'b1), 0 );
$width ( negedge clk &&& (delay_functional_mode == 1'b1), 0 );
$width ( posedge clk &&& (scan_mode == 1'b1), 0 );
$width ( negedge clk &&& (scan_mode == 1'b1), 0 );
$width ( posedge csa_n , 0 ) ;
$width ( negedge csa_n , 0 ) ;
$width ( posedge csb_n , 0 ) ;
$width ( negedge csb_n , 0 ) ;
$width ( posedge dinb , 0 ) ;
$width ( negedge dinb , 0 ) ;
$width ( posedge shift_n , 0 ) ;
$width ( negedge shift_n , 0 ) ;
$width ( posedge sin , 0 ) ;
$width ( negedge sin , 0 ) ;
$period ( posedge clk &&& (delay_functional_mode == 1'b1) , 0 );
$period ( posedge clk &&& (scan_mode == 1'b1) , 0 );
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , posedge addra &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , negedge addra &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , posedge addra &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , negedge addra &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , posedge addrb &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , negedge addrb &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , posedge addrb &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , negedge addrb &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , posedge csa_n &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , negedge csa_n &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , posedge csa_n &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , negedge csa_n &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , posedge csb_n &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , negedge csb_n &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , posedge csb_n &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , negedge csb_n &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , posedge dinb &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( delay_functional_mode == 1'b1) , negedge dinb &&& ( delay_functional_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , posedge dinb &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_capture_mode == 1'b1) , negedge dinb &&& ( scan_capture_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_mode == 1'b1) , posedge shift_n &&& ( scan_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_mode == 1'b1) , negedge shift_n &&& ( scan_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_shift_mode == 1'b1) , posedge sin &&& ( scan_shift_mode == 1'b1 ), 0 , 0 ) ;
$setuphold( posedge clk &&& ( scan_shift_mode == 1'b1) , negedge sin &&& ( scan_shift_mode == 1'b1 ), 0 , 0 ) ;
$setuphold ( posedge clamp_mem, posedge slp_nret_n , 0 , 0 ) ; 
$setuphold ( posedge clamp_mem, negedge slp_nret_n , 0 , 0 ) ; 
$setuphold ( negedge clamp_mem, posedge slp_nret_n , 0 , 0 ) ; 
$setuphold ( negedge clamp_mem, negedge slp_nret_n , 0 , 0 ) ; 
$setuphold ( posedge clamp_mem, posedge slp_ret_n , 0 , 0 ) ; 
$setuphold ( posedge clamp_mem, negedge slp_ret_n , 0 , 0 ) ; 
$setuphold ( negedge clamp_mem, posedge slp_ret_n , 0 , 0 ) ; 
$setuphold ( negedge clamp_mem, negedge slp_ret_n , 0 , 0 ) ; 
endspecify
endmodule 

`endif 


//------> /hd/cad/mentor/2016.9/Mgc_home/pkgs/siflibs/mgc_out_fifo_wait_core_v2001_v9.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_fifo_wait_core_v9 (clk, en, arst, srst, ld, vd, d, lz, vz,  z, sd);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // size of port for elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter integer ph_clk  =  1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en   =  1; // clock enable polarity
    parameter integer ph_arst =  1; // async reset polarity
    parameter integer ph_srst =  1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)

   localparam integer  fifo_b = width * fifo_sz;

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 ld;    // load data
    output                vd;    // fifo full active low
    input     [width-1:0] d;
    output                lz;    // fifo ready to send
    input                 vz;    // dest ready for data
    output    [width-1:0] z;
    output    [sz_width-1:0]      sd; 

    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;
    reg      [fifo_mx:0] stat_pre;
    reg      [fifo_mx:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    wire     [fifo_mx:0] en_l;
    wire     [fifo_mx_over_8:0] en_l_s;

    reg       [width-1:0] buff_nxt;

    reg                   stat_nxt;
    reg                   stat_before;
    reg                   stat_after;
    reg       [fifo_mx:0] en_l_var;

    integer               i;
    genvar                eni;

    wire [32:0]           size_t;
    reg [31:0]            count;
    reg [31:0]            count_t;
    reg [32:0]            n_elem;
    // synopsys translate_off
    reg [31:0]            peak = 32'b0;
    // synopsys translate_on
    wire                  active;

    assign active = ld | vz; // (ld & ~vd) | (vz & ~lz);

    genvar igen;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
      wire [31:0]           delta;
      //  0 :  32'b0      if ld==0 and (vz & stat[fifo_sz-1])==0   
      //               or if ld==1 and (vz & stat[fifo_sz-1])==1
      // +1 :  32'b1      if ld==1 and (vz & stat[fifo_sz-1])==0
      // -1 : {32{1'b1}}  if ld==0 and (vz & stat[fifo_sz-1])==1
      assign delta   =  {{31{(~ld & (vz & stat[fifo_sz-1]))}} , (vz & stat[fifo_sz-1]) ^ ld};
      assign vd = vz | ~stat[0];
      assign lz = ld | stat[fifo_sz-1];
      assign size_t = count + delta;
      assign sd = size_t[sz_width-1:0];
      assign z = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : d;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_before = (i != 0) ? stat[i-1] : 1'b0;
          stat_after = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;
          stat_nxt = stat_after &
                    (stat_before | (stat[i] & (~vz)) | (stat[i] & ld) | (ld & (~vz)));
  
          stat_pre[i] = stat_nxt;
          if (vz & stat_before )
            begin
              buff_nxt[0+:width] = buff[width*(i-1)+:width];
              en_l_var[i] = 1'b1;
            end
          else if (ld & ~((~vz) & stat[i]))
            begin
              buff_nxt = d;
              en_l_var[i] = 1'b1;
            end
          else
            begin
              buff_nxt = d; // Don't care input to disabled flop
              en_l_var[i] = 1'b0;
            end
             
          buff_pre[width*i+:width] = buff_nxt[0+:width];
  
          if ((stat_after == 1'b1) & (stat[i] == 1'b0)) 
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end

        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else 
          count_t = n_elem[31:0];
        count = count_t;
        // synopsys translate_off
        if ( peak < count )
          peak = count;
        // synopsys translate_on
      end

      if (ph_en) begin: PH_EN_HI
        assign en_l_s[fifo_mx_over_8] = en & active;
        for (igen = 0 ; igen < fifo_sz ; igen = igen + 1) begin: NEED_A_LABEL
          assign en_l[igen] = en & en_l_var[igen];
        end
        for (igen = 1 ; igen <= fifo_mx_over_8 ; igen = igen + 1) begin: NEED_A_LABEL2
          assign  en_l_s[igen-1] = en & (stat[igen*8]) & (active);
        end
      end
      else begin: PH_EN_LO
        assign en_l_s[fifo_mx_over_8] = en | ~active;
        for (igen = 0 ; igen < fifo_sz ; igen = igen + 1) begin: NEED_A_LABEL3
          assign en_l[igen] = en | ~en_l_var[igen];
        end
        for (igen = 1 ; igen <= fifo_mx_over_8 ; igen = igen + 1) begin: NEED_A_LABEL2
          assign  en_l_s[igen-1] = en | (~stat[igen*8]) | (~active);
        end
      end

      // Output registers:
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: BUF_GEN
        if (ph_clk==1) begin: POS_BUF
          if (ph_arst==0) begin: LABEL1
            always @(posedge clk or negedge arst)
            if (arst == 1'b0) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
          else begin: LABEL2 // ph_arst==1
            always @(posedge clk or posedge arst)
            if (arst == 1'b1) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
        end
        else begin: NEG_BUF
          if (ph_arst==0) begin: LABEL3
            always @(negedge clk or negedge arst)
            if (arst == 1'b0) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
          else begin: LABEL4 // ph_arst==1
            always @(negedge clk or posedge arst)
            if (arst == 1'b1) begin
              stat[eni] <= 1'b0;
            end
            else if (srst == ph_srst) begin
              stat[eni] <= 1'b0;
            end
            else if (en_l_s[eni/8] == ph_en) begin
              stat[eni] <= stat_pre[eni];
            end
          end
        end
      end

      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: STATGEN2
        if (ph_clk==1) begin: POS_STAT
          if (ph_arst==0) begin: LABEL5
            always @(posedge clk or negedge arst)
            if (arst == 1'b0) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
          else begin: LABEL6 // ph_arst==1
            always @(posedge clk or posedge arst)
            if (arst == 1'b1) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
        end
        else begin: NEG_STAT // ph_clk==0
          if (ph_arst==0) begin: LABEL7
            always @(negedge clk or negedge arst)
            if (arst == 1'b0) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
          else begin: LABEL8 // ph_arst==1
            always @(negedge clk or posedge arst)
            if (arst == 1'b1) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (srst == ph_srst) begin
              buff[width*eni+:width] <= {width{1'b0}};
            end
            else if (en_l[eni] == ph_en) begin
              buff[width*eni+:width] <= buff_pre[width*eni+:width];
            end
          end
        end
      end
    end
    else
    begin: FEED_THRU
      assign vd = vz;
      assign lz = ld;
      assign z = d;
      assign sd = ld & ~vz;
    end
    endgenerate

endmodule



//------> /hd/cad/mentor/2016.9/Mgc_home/pkgs/siflibs/mgc_pipe_v2001_v10.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


/*
 *
 *             _______________________________________________
 * WRITER    |                                               |          READER
 *           |           MGC_PIPE                            |
 *           |           __________________________          |
 *        --<| vdout  --<| vd ---------------  vz<|-----ldin<|---
 *           |           |      FIFO              |          |
 *        ---|>ldout  ---|>ld ---------------- lz |> ---vdin |>--
 *        ---|>dout -----|>d  ---------------- dz |> ----din |>--
 *           |           |________________________|          |
 *           |_______________________________________________|
 *
 *    vdout - can be considered as a notFULL signal
 *    vdin  - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from ldout & !vdout
 *    read_stall  - an internal debug signal formed from ldin & !vdin
 *
 */
// two clock pipe
module mgc_pipe_v10 (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, sd);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter integer log2_sz = 3; // log2(fifo_sz)
    parameter integer ph_clk  = 1;  // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en   = 1;  // clock enable polarity
    parameter integer ph_arst = 1;  // async reset polarity
    parameter integer ph_srst = 1;  // sync reset polarity

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output [sz_width-1:0]      sd;

    // synopsys translate_off
    wire               write_stall;
    wire               read_stall;
    assign write_stall = ldout & !vdout;
    assign read_stall = ldin & !vdin;
    // synopsys translate_on

    mgc_out_fifo_wait_core_v9
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz)
    )
    FIFO
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (vdin),
        .vz      (ldin),
        .z       (din),
        .sd      (sd)
    );

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/263344 Production Release
//  HLS Date:       Sun Jul  3 19:13:39 PDT 2016
// 
//  Generated by:   xuany@kiwi
//  Generated date: Wed Mar 28 17:40:27 2018
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    double_buffeoFsRV17_cns_bctl
// ------------------------------------------------------------------


module double_buffeoFsRV17_cns_bctl (
  clk, rst, dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_17_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_17_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_17_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_17_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_17_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_17_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_17_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_17_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_17_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_17_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_17_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_17_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_17_cns_S0, shr_mem_17_cns_R0, shr_mem_17_cns_S1, shr_mem_17_cns_R1,
      shr_mem_17_cns_addra_shi0, shr_mem_17_cns_addra_shi1, shr_mem_17_cns_addrb_shi0,
      shr_mem_17_cns_addrb_shi1, shr_mem_17_cns_csa_n_shi0, shr_mem_17_cns_csa_n_shi1,
      shr_mem_17_cns_csb_n_shi0, shr_mem_17_cns_csb_n_shi1, shr_mem_17_cns_dinb_shi0,
      shr_mem_17_cns_dinb_shi1, shr_mem_17_cns_douta_sho0, shr_mem_17_cns_douta_sho1,
      shr_mem_17_cns_S1_pff, din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_17_cns_S0_pff
);
  input clk;
  input rst;
  input dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_17_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_17_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_17_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_17_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_17_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_17_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_17_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_17_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_17_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_17_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_17_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_17_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_17_cns_S0;
  input shr_mem_17_cns_R0;
  output shr_mem_17_cns_S1;
  input shr_mem_17_cns_R1;
  output [6:0] shr_mem_17_cns_addra_shi0;
  output [6:0] shr_mem_17_cns_addra_shi1;
  output [6:0] shr_mem_17_cns_addrb_shi0;
  output [6:0] shr_mem_17_cns_addrb_shi1;
  output shr_mem_17_cns_csa_n_shi0;
  output shr_mem_17_cns_csa_n_shi1;
  output shr_mem_17_cns_csb_n_shi0;
  output shr_mem_17_cns_csb_n_shi1;
  output [63:0] shr_mem_17_cns_dinb_shi0;
  output [63:0] shr_mem_17_cns_dinb_shi1;
  input [63:0] shr_mem_17_cns_douta_sho0;
  input [63:0] shr_mem_17_cns_douta_sho1;
  output shr_mem_17_cns_S1_pff;
  input din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_17_cns_S0_pff;


  // Interconnect Declarations
  reg dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_17_cns_PC0;
  reg shr_mem_17_cns_ppidx;
  reg [1:0] shr_mem_17_cns_ppown;
  wire shr_mem_17_cns_PC1;
  reg shr_mem_17_cns_ppidx_1;
  reg [1:0] shr_mem_17_cns_ppown_1;
  wire [6:0] shr_mem_17_shr_mem_17_mux_3_cse_pff;
  wire shr_mem_17_and_3_cse_pff;
  wire [1:0] shr_mem_17_acc_1_rmff;
  wire [3:0] nl_shr_mem_17_acc_1_rmff;
  wire shr_mem_17_xor_1_rmff;
  wire shr_mem_17_shr_mem_17_or_cse_pff;
  wire [1:0] shr_mem_17_acc_rmff;
  wire [3:0] nl_shr_mem_17_acc_rmff;
  wire shr_mem_17_xor_rmff;
  wire [6:0] shr_mem_17_shr_mem_17_mux_2_cse_pff;
  wire shr_mem_17_and_5_cse_pff;
  wire shr_mem_17_shr_mem_17_or_1_cse_pff;

  wire[0:0] shr_mem_17_mux_6_nl;
  wire[0:0] shr_mem_17_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_17_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_17_cns_R0;
  assign din_17_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_17_cns_R1;
  assign shr_mem_17_xor_rmff = shr_mem_17_cns_ppidx ^ shr_mem_17_cns_PC0;
  assign nl_shr_mem_17_acc_rmff = shr_mem_17_cns_ppown + conv_u2u_1_2(shr_mem_17_cns_PC0)
      + conv_s2u_1_2(shr_mem_17_cns_PC1);
  assign shr_mem_17_acc_rmff = nl_shr_mem_17_acc_rmff[1:0];
  assign shr_mem_17_cns_PC0 = shr_mem_17_cns_S0 & dout_17_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_17_xor_1_rmff = shr_mem_17_cns_ppidx_1 ^ shr_mem_17_cns_PC1;
  assign nl_shr_mem_17_acc_1_rmff = shr_mem_17_cns_ppown_1 + conv_u2u_1_2(shr_mem_17_cns_PC1)
      + conv_s2u_1_2(shr_mem_17_cns_PC0);
  assign shr_mem_17_acc_1_rmff = nl_shr_mem_17_acc_1_rmff[1:0];
  assign shr_mem_17_cns_PC1 = shr_mem_17_cns_S1 & din_17_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_17_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_17_cns_douta_sho0,
      shr_mem_17_cns_douta_sho1, shr_mem_17_cns_ppidx);
  assign din_17_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_17_cns_douta_sho0,
      shr_mem_17_cns_douta_sho1, shr_mem_17_cns_ppidx_1);
  assign shr_mem_17_cns_addra_shi0 = shr_mem_17_shr_mem_17_mux_3_cse_pff;
  assign shr_mem_17_cns_S1 = (shr_mem_17_cns_ppown_1!=2'b00);
  assign shr_mem_17_cns_S1_pff = (shr_mem_17_acc_1_rmff!=2'b00);
  assign shr_mem_17_and_3_cse_pff = shr_mem_17_cns_S1_pff & (~ shr_mem_17_xor_1_rmff);
  assign shr_mem_17_shr_mem_17_mux_3_cse_pff = MUX_v_7_2_2(dout_17_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_17_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_17_and_3_cse_pff);
  assign shr_mem_17_cns_addrb_shi0 = shr_mem_17_shr_mem_17_mux_3_cse_pff;
  assign shr_mem_17_cns_csa_n_shi0 = shr_mem_17_shr_mem_17_or_cse_pff;
  assign din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff =
      din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff =
      dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_17_cns_S0 = ~((shr_mem_17_cns_ppown==2'b10));
  assign shr_mem_17_cns_S0_pff = ~((shr_mem_17_acc_rmff==2'b10));
  assign shr_mem_17_mux_6_nl = MUX_s_1_2_2(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_17_and_3_cse_pff);
  assign shr_mem_17_shr_mem_17_or_cse_pff = (shr_mem_17_mux_6_nl) | (~((shr_mem_17_cns_S0_pff
      & (~ shr_mem_17_xor_rmff)) | shr_mem_17_and_3_cse_pff));
  assign shr_mem_17_cns_csb_n_shi0 = shr_mem_17_shr_mem_17_or_cse_pff;
  assign shr_mem_17_cns_dinb_shi0 = MUX_v_64_2_2(dout_17_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_17_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_17_and_3_cse_pff);
  assign shr_mem_17_cns_addra_shi1 = shr_mem_17_shr_mem_17_mux_2_cse_pff;
  assign shr_mem_17_and_5_cse_pff = shr_mem_17_cns_S1_pff & shr_mem_17_xor_1_rmff;
  assign shr_mem_17_shr_mem_17_mux_2_cse_pff = MUX_v_7_2_2(dout_17_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_17_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_17_and_5_cse_pff);
  assign shr_mem_17_cns_addrb_shi1 = shr_mem_17_shr_mem_17_mux_2_cse_pff;
  assign shr_mem_17_cns_csa_n_shi1 = shr_mem_17_shr_mem_17_or_1_cse_pff;
  assign shr_mem_17_mux_7_nl = MUX_s_1_2_2(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_17_and_5_cse_pff);
  assign shr_mem_17_shr_mem_17_or_1_cse_pff = (shr_mem_17_mux_7_nl) | (~((shr_mem_17_cns_S0_pff
      & shr_mem_17_xor_rmff) | shr_mem_17_and_5_cse_pff));
  assign shr_mem_17_cns_csb_n_shi1 = shr_mem_17_shr_mem_17_or_1_cse_pff;
  assign shr_mem_17_cns_dinb_shi1 = MUX_v_64_2_2(dout_17_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_17_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_17_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_17_cns_ppidx <= 1'b0;
      shr_mem_17_cns_ppown <= 2'b0;
      shr_mem_17_cns_ppidx_1 <= 1'b0;
      shr_mem_17_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_17_cns_ppidx <= shr_mem_17_xor_rmff;
      shr_mem_17_cns_ppown <= shr_mem_17_acc_rmff;
      shr_mem_17_cns_ppidx_1 <= shr_mem_17_xor_1_rmff;
      shr_mem_17_cns_ppown_1 <= shr_mem_17_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeoFsRV16_cns_bctl
// ------------------------------------------------------------------


module double_buffeoFsRV16_cns_bctl (
  clk, rst, dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_16_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_16_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_16_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_16_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_16_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_16_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_16_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_16_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_16_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_16_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_16_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_16_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_16_cns_S0, shr_mem_16_cns_R0, shr_mem_16_cns_S1, shr_mem_16_cns_R1,
      shr_mem_16_cns_addra_shi0, shr_mem_16_cns_addra_shi1, shr_mem_16_cns_addrb_shi0,
      shr_mem_16_cns_addrb_shi1, shr_mem_16_cns_csa_n_shi0, shr_mem_16_cns_csa_n_shi1,
      shr_mem_16_cns_csb_n_shi0, shr_mem_16_cns_csb_n_shi1, shr_mem_16_cns_dinb_shi0,
      shr_mem_16_cns_dinb_shi1, shr_mem_16_cns_douta_sho0, shr_mem_16_cns_douta_sho1,
      shr_mem_16_cns_S1_pff, din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_16_cns_S0_pff
);
  input clk;
  input rst;
  input dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_16_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_16_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_16_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_16_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_16_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_16_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_16_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_16_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_16_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_16_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_16_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_16_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_16_cns_S0;
  input shr_mem_16_cns_R0;
  output shr_mem_16_cns_S1;
  input shr_mem_16_cns_R1;
  output [6:0] shr_mem_16_cns_addra_shi0;
  output [6:0] shr_mem_16_cns_addra_shi1;
  output [6:0] shr_mem_16_cns_addrb_shi0;
  output [6:0] shr_mem_16_cns_addrb_shi1;
  output shr_mem_16_cns_csa_n_shi0;
  output shr_mem_16_cns_csa_n_shi1;
  output shr_mem_16_cns_csb_n_shi0;
  output shr_mem_16_cns_csb_n_shi1;
  output [63:0] shr_mem_16_cns_dinb_shi0;
  output [63:0] shr_mem_16_cns_dinb_shi1;
  input [63:0] shr_mem_16_cns_douta_sho0;
  input [63:0] shr_mem_16_cns_douta_sho1;
  output shr_mem_16_cns_S1_pff;
  input din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_16_cns_S0_pff;


  // Interconnect Declarations
  reg dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_16_cns_PC0;
  reg shr_mem_16_cns_ppidx;
  reg [1:0] shr_mem_16_cns_ppown;
  wire shr_mem_16_cns_PC1;
  reg shr_mem_16_cns_ppidx_1;
  reg [1:0] shr_mem_16_cns_ppown_1;
  wire [6:0] shr_mem_16_shr_mem_16_mux_3_cse_pff;
  wire shr_mem_16_and_3_cse_pff;
  wire [1:0] shr_mem_16_acc_1_rmff;
  wire [3:0] nl_shr_mem_16_acc_1_rmff;
  wire shr_mem_16_xor_1_rmff;
  wire shr_mem_16_shr_mem_16_or_cse_pff;
  wire [1:0] shr_mem_16_acc_rmff;
  wire [3:0] nl_shr_mem_16_acc_rmff;
  wire shr_mem_16_xor_rmff;
  wire [6:0] shr_mem_16_shr_mem_16_mux_2_cse_pff;
  wire shr_mem_16_and_5_cse_pff;
  wire shr_mem_16_shr_mem_16_or_1_cse_pff;

  wire[0:0] shr_mem_16_mux_6_nl;
  wire[0:0] shr_mem_16_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_16_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_16_cns_R0;
  assign din_16_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_16_cns_R1;
  assign shr_mem_16_xor_rmff = shr_mem_16_cns_ppidx ^ shr_mem_16_cns_PC0;
  assign nl_shr_mem_16_acc_rmff = shr_mem_16_cns_ppown + conv_u2u_1_2(shr_mem_16_cns_PC0)
      + conv_s2u_1_2(shr_mem_16_cns_PC1);
  assign shr_mem_16_acc_rmff = nl_shr_mem_16_acc_rmff[1:0];
  assign shr_mem_16_cns_PC0 = shr_mem_16_cns_S0 & dout_16_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_16_xor_1_rmff = shr_mem_16_cns_ppidx_1 ^ shr_mem_16_cns_PC1;
  assign nl_shr_mem_16_acc_1_rmff = shr_mem_16_cns_ppown_1 + conv_u2u_1_2(shr_mem_16_cns_PC1)
      + conv_s2u_1_2(shr_mem_16_cns_PC0);
  assign shr_mem_16_acc_1_rmff = nl_shr_mem_16_acc_1_rmff[1:0];
  assign shr_mem_16_cns_PC1 = shr_mem_16_cns_S1 & din_16_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_16_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_16_cns_douta_sho0,
      shr_mem_16_cns_douta_sho1, shr_mem_16_cns_ppidx);
  assign din_16_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_16_cns_douta_sho0,
      shr_mem_16_cns_douta_sho1, shr_mem_16_cns_ppidx_1);
  assign shr_mem_16_cns_addra_shi0 = shr_mem_16_shr_mem_16_mux_3_cse_pff;
  assign shr_mem_16_cns_S1 = (shr_mem_16_cns_ppown_1!=2'b00);
  assign shr_mem_16_cns_S1_pff = (shr_mem_16_acc_1_rmff!=2'b00);
  assign shr_mem_16_and_3_cse_pff = shr_mem_16_cns_S1_pff & (~ shr_mem_16_xor_1_rmff);
  assign shr_mem_16_shr_mem_16_mux_3_cse_pff = MUX_v_7_2_2(dout_16_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_16_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_16_and_3_cse_pff);
  assign shr_mem_16_cns_addrb_shi0 = shr_mem_16_shr_mem_16_mux_3_cse_pff;
  assign shr_mem_16_cns_csa_n_shi0 = shr_mem_16_shr_mem_16_or_cse_pff;
  assign din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff =
      din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff =
      dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_16_cns_S0 = ~((shr_mem_16_cns_ppown==2'b10));
  assign shr_mem_16_cns_S0_pff = ~((shr_mem_16_acc_rmff==2'b10));
  assign shr_mem_16_mux_6_nl = MUX_s_1_2_2(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_16_and_3_cse_pff);
  assign shr_mem_16_shr_mem_16_or_cse_pff = (shr_mem_16_mux_6_nl) | (~((shr_mem_16_cns_S0_pff
      & (~ shr_mem_16_xor_rmff)) | shr_mem_16_and_3_cse_pff));
  assign shr_mem_16_cns_csb_n_shi0 = shr_mem_16_shr_mem_16_or_cse_pff;
  assign shr_mem_16_cns_dinb_shi0 = MUX_v_64_2_2(dout_16_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_16_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_16_and_3_cse_pff);
  assign shr_mem_16_cns_addra_shi1 = shr_mem_16_shr_mem_16_mux_2_cse_pff;
  assign shr_mem_16_and_5_cse_pff = shr_mem_16_cns_S1_pff & shr_mem_16_xor_1_rmff;
  assign shr_mem_16_shr_mem_16_mux_2_cse_pff = MUX_v_7_2_2(dout_16_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_16_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_16_and_5_cse_pff);
  assign shr_mem_16_cns_addrb_shi1 = shr_mem_16_shr_mem_16_mux_2_cse_pff;
  assign shr_mem_16_cns_csa_n_shi1 = shr_mem_16_shr_mem_16_or_1_cse_pff;
  assign shr_mem_16_mux_7_nl = MUX_s_1_2_2(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_16_and_5_cse_pff);
  assign shr_mem_16_shr_mem_16_or_1_cse_pff = (shr_mem_16_mux_7_nl) | (~((shr_mem_16_cns_S0_pff
      & shr_mem_16_xor_rmff) | shr_mem_16_and_5_cse_pff));
  assign shr_mem_16_cns_csb_n_shi1 = shr_mem_16_shr_mem_16_or_1_cse_pff;
  assign shr_mem_16_cns_dinb_shi1 = MUX_v_64_2_2(dout_16_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_16_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_16_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_16_cns_ppidx <= 1'b0;
      shr_mem_16_cns_ppown <= 2'b0;
      shr_mem_16_cns_ppidx_1 <= 1'b0;
      shr_mem_16_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_16_cns_ppidx <= shr_mem_16_xor_rmff;
      shr_mem_16_cns_ppown <= shr_mem_16_acc_rmff;
      shr_mem_16_cns_ppidx_1 <= shr_mem_16_xor_1_rmff;
      shr_mem_16_cns_ppown_1 <= shr_mem_16_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeoFsRV15_cns_bctl
// ------------------------------------------------------------------


module double_buffeoFsRV15_cns_bctl (
  clk, rst, dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_15_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_15_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_15_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_15_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_15_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_15_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_15_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_15_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_15_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_15_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_15_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_15_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_15_cns_S0, shr_mem_15_cns_R0, shr_mem_15_cns_S1, shr_mem_15_cns_R1,
      shr_mem_15_cns_addra_shi0, shr_mem_15_cns_addra_shi1, shr_mem_15_cns_addrb_shi0,
      shr_mem_15_cns_addrb_shi1, shr_mem_15_cns_csa_n_shi0, shr_mem_15_cns_csa_n_shi1,
      shr_mem_15_cns_csb_n_shi0, shr_mem_15_cns_csb_n_shi1, shr_mem_15_cns_dinb_shi0,
      shr_mem_15_cns_dinb_shi1, shr_mem_15_cns_douta_sho0, shr_mem_15_cns_douta_sho1,
      shr_mem_15_cns_S1_pff, din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_15_cns_S0_pff
);
  input clk;
  input rst;
  input dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_15_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_15_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_15_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_15_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_15_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_15_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_15_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_15_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_15_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_15_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_15_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_15_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_15_cns_S0;
  input shr_mem_15_cns_R0;
  output shr_mem_15_cns_S1;
  input shr_mem_15_cns_R1;
  output [6:0] shr_mem_15_cns_addra_shi0;
  output [6:0] shr_mem_15_cns_addra_shi1;
  output [6:0] shr_mem_15_cns_addrb_shi0;
  output [6:0] shr_mem_15_cns_addrb_shi1;
  output shr_mem_15_cns_csa_n_shi0;
  output shr_mem_15_cns_csa_n_shi1;
  output shr_mem_15_cns_csb_n_shi0;
  output shr_mem_15_cns_csb_n_shi1;
  output [63:0] shr_mem_15_cns_dinb_shi0;
  output [63:0] shr_mem_15_cns_dinb_shi1;
  input [63:0] shr_mem_15_cns_douta_sho0;
  input [63:0] shr_mem_15_cns_douta_sho1;
  output shr_mem_15_cns_S1_pff;
  input din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_15_cns_S0_pff;


  // Interconnect Declarations
  reg dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_15_cns_PC0;
  reg shr_mem_15_cns_ppidx;
  reg [1:0] shr_mem_15_cns_ppown;
  wire shr_mem_15_cns_PC1;
  reg shr_mem_15_cns_ppidx_1;
  reg [1:0] shr_mem_15_cns_ppown_1;
  wire [6:0] shr_mem_15_shr_mem_15_mux_3_cse_pff;
  wire shr_mem_15_and_3_cse_pff;
  wire [1:0] shr_mem_15_acc_1_rmff;
  wire [3:0] nl_shr_mem_15_acc_1_rmff;
  wire shr_mem_15_xor_1_rmff;
  wire shr_mem_15_shr_mem_15_or_cse_pff;
  wire [1:0] shr_mem_15_acc_rmff;
  wire [3:0] nl_shr_mem_15_acc_rmff;
  wire shr_mem_15_xor_rmff;
  wire [6:0] shr_mem_15_shr_mem_15_mux_2_cse_pff;
  wire shr_mem_15_and_5_cse_pff;
  wire shr_mem_15_shr_mem_15_or_1_cse_pff;

  wire[0:0] shr_mem_15_mux_6_nl;
  wire[0:0] shr_mem_15_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_15_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_15_cns_R0;
  assign din_15_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_15_cns_R1;
  assign shr_mem_15_xor_rmff = shr_mem_15_cns_ppidx ^ shr_mem_15_cns_PC0;
  assign nl_shr_mem_15_acc_rmff = shr_mem_15_cns_ppown + conv_u2u_1_2(shr_mem_15_cns_PC0)
      + conv_s2u_1_2(shr_mem_15_cns_PC1);
  assign shr_mem_15_acc_rmff = nl_shr_mem_15_acc_rmff[1:0];
  assign shr_mem_15_cns_PC0 = shr_mem_15_cns_S0 & dout_15_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_15_xor_1_rmff = shr_mem_15_cns_ppidx_1 ^ shr_mem_15_cns_PC1;
  assign nl_shr_mem_15_acc_1_rmff = shr_mem_15_cns_ppown_1 + conv_u2u_1_2(shr_mem_15_cns_PC1)
      + conv_s2u_1_2(shr_mem_15_cns_PC0);
  assign shr_mem_15_acc_1_rmff = nl_shr_mem_15_acc_1_rmff[1:0];
  assign shr_mem_15_cns_PC1 = shr_mem_15_cns_S1 & din_15_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_15_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_15_cns_douta_sho0,
      shr_mem_15_cns_douta_sho1, shr_mem_15_cns_ppidx);
  assign din_15_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_15_cns_douta_sho0,
      shr_mem_15_cns_douta_sho1, shr_mem_15_cns_ppidx_1);
  assign shr_mem_15_cns_addra_shi0 = shr_mem_15_shr_mem_15_mux_3_cse_pff;
  assign shr_mem_15_cns_S1 = (shr_mem_15_cns_ppown_1!=2'b00);
  assign shr_mem_15_cns_S1_pff = (shr_mem_15_acc_1_rmff!=2'b00);
  assign shr_mem_15_and_3_cse_pff = shr_mem_15_cns_S1_pff & (~ shr_mem_15_xor_1_rmff);
  assign shr_mem_15_shr_mem_15_mux_3_cse_pff = MUX_v_7_2_2(dout_15_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_15_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_15_and_3_cse_pff);
  assign shr_mem_15_cns_addrb_shi0 = shr_mem_15_shr_mem_15_mux_3_cse_pff;
  assign shr_mem_15_cns_csa_n_shi0 = shr_mem_15_shr_mem_15_or_cse_pff;
  assign din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff =
      din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff =
      dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_15_cns_S0 = ~((shr_mem_15_cns_ppown==2'b10));
  assign shr_mem_15_cns_S0_pff = ~((shr_mem_15_acc_rmff==2'b10));
  assign shr_mem_15_mux_6_nl = MUX_s_1_2_2(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_15_and_3_cse_pff);
  assign shr_mem_15_shr_mem_15_or_cse_pff = (shr_mem_15_mux_6_nl) | (~((shr_mem_15_cns_S0_pff
      & (~ shr_mem_15_xor_rmff)) | shr_mem_15_and_3_cse_pff));
  assign shr_mem_15_cns_csb_n_shi0 = shr_mem_15_shr_mem_15_or_cse_pff;
  assign shr_mem_15_cns_dinb_shi0 = MUX_v_64_2_2(dout_15_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_15_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_15_and_3_cse_pff);
  assign shr_mem_15_cns_addra_shi1 = shr_mem_15_shr_mem_15_mux_2_cse_pff;
  assign shr_mem_15_and_5_cse_pff = shr_mem_15_cns_S1_pff & shr_mem_15_xor_1_rmff;
  assign shr_mem_15_shr_mem_15_mux_2_cse_pff = MUX_v_7_2_2(dout_15_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_15_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_15_and_5_cse_pff);
  assign shr_mem_15_cns_addrb_shi1 = shr_mem_15_shr_mem_15_mux_2_cse_pff;
  assign shr_mem_15_cns_csa_n_shi1 = shr_mem_15_shr_mem_15_or_1_cse_pff;
  assign shr_mem_15_mux_7_nl = MUX_s_1_2_2(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_15_and_5_cse_pff);
  assign shr_mem_15_shr_mem_15_or_1_cse_pff = (shr_mem_15_mux_7_nl) | (~((shr_mem_15_cns_S0_pff
      & shr_mem_15_xor_rmff) | shr_mem_15_and_5_cse_pff));
  assign shr_mem_15_cns_csb_n_shi1 = shr_mem_15_shr_mem_15_or_1_cse_pff;
  assign shr_mem_15_cns_dinb_shi1 = MUX_v_64_2_2(dout_15_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_15_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_15_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_15_cns_ppidx <= 1'b0;
      shr_mem_15_cns_ppown <= 2'b0;
      shr_mem_15_cns_ppidx_1 <= 1'b0;
      shr_mem_15_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_15_cns_ppidx <= shr_mem_15_xor_rmff;
      shr_mem_15_cns_ppown <= shr_mem_15_acc_rmff;
      shr_mem_15_cns_ppidx_1 <= shr_mem_15_xor_1_rmff;
      shr_mem_15_cns_ppown_1 <= shr_mem_15_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeoFsRV14_cns_bctl
// ------------------------------------------------------------------


module double_buffeoFsRV14_cns_bctl (
  clk, rst, dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_14_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_14_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_14_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_14_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_14_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_14_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_14_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_14_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_14_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_14_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_14_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_14_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_14_cns_S0, shr_mem_14_cns_R0, shr_mem_14_cns_S1, shr_mem_14_cns_R1,
      shr_mem_14_cns_addra_shi0, shr_mem_14_cns_addra_shi1, shr_mem_14_cns_addrb_shi0,
      shr_mem_14_cns_addrb_shi1, shr_mem_14_cns_csa_n_shi0, shr_mem_14_cns_csa_n_shi1,
      shr_mem_14_cns_csb_n_shi0, shr_mem_14_cns_csb_n_shi1, shr_mem_14_cns_dinb_shi0,
      shr_mem_14_cns_dinb_shi1, shr_mem_14_cns_douta_sho0, shr_mem_14_cns_douta_sho1,
      shr_mem_14_cns_S1_pff, din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_14_cns_S0_pff
);
  input clk;
  input rst;
  input dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_14_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_14_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_14_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_14_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_14_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_14_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_14_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_14_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_14_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_14_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_14_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_14_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_14_cns_S0;
  input shr_mem_14_cns_R0;
  output shr_mem_14_cns_S1;
  input shr_mem_14_cns_R1;
  output [6:0] shr_mem_14_cns_addra_shi0;
  output [6:0] shr_mem_14_cns_addra_shi1;
  output [6:0] shr_mem_14_cns_addrb_shi0;
  output [6:0] shr_mem_14_cns_addrb_shi1;
  output shr_mem_14_cns_csa_n_shi0;
  output shr_mem_14_cns_csa_n_shi1;
  output shr_mem_14_cns_csb_n_shi0;
  output shr_mem_14_cns_csb_n_shi1;
  output [63:0] shr_mem_14_cns_dinb_shi0;
  output [63:0] shr_mem_14_cns_dinb_shi1;
  input [63:0] shr_mem_14_cns_douta_sho0;
  input [63:0] shr_mem_14_cns_douta_sho1;
  output shr_mem_14_cns_S1_pff;
  input din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_14_cns_S0_pff;


  // Interconnect Declarations
  reg dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_14_cns_PC0;
  reg shr_mem_14_cns_ppidx;
  reg [1:0] shr_mem_14_cns_ppown;
  wire shr_mem_14_cns_PC1;
  reg shr_mem_14_cns_ppidx_1;
  reg [1:0] shr_mem_14_cns_ppown_1;
  wire [6:0] shr_mem_14_shr_mem_14_mux_3_cse_pff;
  wire shr_mem_14_and_3_cse_pff;
  wire [1:0] shr_mem_14_acc_1_rmff;
  wire [3:0] nl_shr_mem_14_acc_1_rmff;
  wire shr_mem_14_xor_1_rmff;
  wire shr_mem_14_shr_mem_14_or_cse_pff;
  wire [1:0] shr_mem_14_acc_rmff;
  wire [3:0] nl_shr_mem_14_acc_rmff;
  wire shr_mem_14_xor_rmff;
  wire [6:0] shr_mem_14_shr_mem_14_mux_2_cse_pff;
  wire shr_mem_14_and_5_cse_pff;
  wire shr_mem_14_shr_mem_14_or_1_cse_pff;

  wire[0:0] shr_mem_14_mux_6_nl;
  wire[0:0] shr_mem_14_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_14_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_14_cns_R0;
  assign din_14_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_14_cns_R1;
  assign shr_mem_14_xor_rmff = shr_mem_14_cns_ppidx ^ shr_mem_14_cns_PC0;
  assign nl_shr_mem_14_acc_rmff = shr_mem_14_cns_ppown + conv_u2u_1_2(shr_mem_14_cns_PC0)
      + conv_s2u_1_2(shr_mem_14_cns_PC1);
  assign shr_mem_14_acc_rmff = nl_shr_mem_14_acc_rmff[1:0];
  assign shr_mem_14_cns_PC0 = shr_mem_14_cns_S0 & dout_14_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_14_xor_1_rmff = shr_mem_14_cns_ppidx_1 ^ shr_mem_14_cns_PC1;
  assign nl_shr_mem_14_acc_1_rmff = shr_mem_14_cns_ppown_1 + conv_u2u_1_2(shr_mem_14_cns_PC1)
      + conv_s2u_1_2(shr_mem_14_cns_PC0);
  assign shr_mem_14_acc_1_rmff = nl_shr_mem_14_acc_1_rmff[1:0];
  assign shr_mem_14_cns_PC1 = shr_mem_14_cns_S1 & din_14_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_14_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_14_cns_douta_sho0,
      shr_mem_14_cns_douta_sho1, shr_mem_14_cns_ppidx);
  assign din_14_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_14_cns_douta_sho0,
      shr_mem_14_cns_douta_sho1, shr_mem_14_cns_ppidx_1);
  assign shr_mem_14_cns_addra_shi0 = shr_mem_14_shr_mem_14_mux_3_cse_pff;
  assign shr_mem_14_cns_S1 = (shr_mem_14_cns_ppown_1!=2'b00);
  assign shr_mem_14_cns_S1_pff = (shr_mem_14_acc_1_rmff!=2'b00);
  assign shr_mem_14_and_3_cse_pff = shr_mem_14_cns_S1_pff & (~ shr_mem_14_xor_1_rmff);
  assign shr_mem_14_shr_mem_14_mux_3_cse_pff = MUX_v_7_2_2(dout_14_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_14_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_14_and_3_cse_pff);
  assign shr_mem_14_cns_addrb_shi0 = shr_mem_14_shr_mem_14_mux_3_cse_pff;
  assign shr_mem_14_cns_csa_n_shi0 = shr_mem_14_shr_mem_14_or_cse_pff;
  assign din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff =
      din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff =
      dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_14_cns_S0 = ~((shr_mem_14_cns_ppown==2'b10));
  assign shr_mem_14_cns_S0_pff = ~((shr_mem_14_acc_rmff==2'b10));
  assign shr_mem_14_mux_6_nl = MUX_s_1_2_2(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_14_and_3_cse_pff);
  assign shr_mem_14_shr_mem_14_or_cse_pff = (shr_mem_14_mux_6_nl) | (~((shr_mem_14_cns_S0_pff
      & (~ shr_mem_14_xor_rmff)) | shr_mem_14_and_3_cse_pff));
  assign shr_mem_14_cns_csb_n_shi0 = shr_mem_14_shr_mem_14_or_cse_pff;
  assign shr_mem_14_cns_dinb_shi0 = MUX_v_64_2_2(dout_14_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_14_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_14_and_3_cse_pff);
  assign shr_mem_14_cns_addra_shi1 = shr_mem_14_shr_mem_14_mux_2_cse_pff;
  assign shr_mem_14_and_5_cse_pff = shr_mem_14_cns_S1_pff & shr_mem_14_xor_1_rmff;
  assign shr_mem_14_shr_mem_14_mux_2_cse_pff = MUX_v_7_2_2(dout_14_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_14_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_14_and_5_cse_pff);
  assign shr_mem_14_cns_addrb_shi1 = shr_mem_14_shr_mem_14_mux_2_cse_pff;
  assign shr_mem_14_cns_csa_n_shi1 = shr_mem_14_shr_mem_14_or_1_cse_pff;
  assign shr_mem_14_mux_7_nl = MUX_s_1_2_2(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_14_and_5_cse_pff);
  assign shr_mem_14_shr_mem_14_or_1_cse_pff = (shr_mem_14_mux_7_nl) | (~((shr_mem_14_cns_S0_pff
      & shr_mem_14_xor_rmff) | shr_mem_14_and_5_cse_pff));
  assign shr_mem_14_cns_csb_n_shi1 = shr_mem_14_shr_mem_14_or_1_cse_pff;
  assign shr_mem_14_cns_dinb_shi1 = MUX_v_64_2_2(dout_14_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_14_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_14_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_14_cns_ppidx <= 1'b0;
      shr_mem_14_cns_ppown <= 2'b0;
      shr_mem_14_cns_ppidx_1 <= 1'b0;
      shr_mem_14_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_14_cns_ppidx <= shr_mem_14_xor_rmff;
      shr_mem_14_cns_ppown <= shr_mem_14_acc_rmff;
      shr_mem_14_cns_ppidx_1 <= shr_mem_14_xor_1_rmff;
      shr_mem_14_cns_ppown_1 <= shr_mem_14_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeoFsRV13_cns_bctl
// ------------------------------------------------------------------


module double_buffeoFsRV13_cns_bctl (
  clk, rst, dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_13_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_13_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_13_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_13_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_13_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_13_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_13_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_13_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_13_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_13_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_13_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_13_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_13_cns_S0, shr_mem_13_cns_R0, shr_mem_13_cns_S1, shr_mem_13_cns_R1,
      shr_mem_13_cns_addra_shi0, shr_mem_13_cns_addra_shi1, shr_mem_13_cns_addrb_shi0,
      shr_mem_13_cns_addrb_shi1, shr_mem_13_cns_csa_n_shi0, shr_mem_13_cns_csa_n_shi1,
      shr_mem_13_cns_csb_n_shi0, shr_mem_13_cns_csb_n_shi1, shr_mem_13_cns_dinb_shi0,
      shr_mem_13_cns_dinb_shi1, shr_mem_13_cns_douta_sho0, shr_mem_13_cns_douta_sho1,
      shr_mem_13_cns_S1_pff, din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_13_cns_S0_pff
);
  input clk;
  input rst;
  input dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_13_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_13_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_13_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_13_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_13_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_13_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_13_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_13_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_13_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_13_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_13_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_13_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_13_cns_S0;
  input shr_mem_13_cns_R0;
  output shr_mem_13_cns_S1;
  input shr_mem_13_cns_R1;
  output [6:0] shr_mem_13_cns_addra_shi0;
  output [6:0] shr_mem_13_cns_addra_shi1;
  output [6:0] shr_mem_13_cns_addrb_shi0;
  output [6:0] shr_mem_13_cns_addrb_shi1;
  output shr_mem_13_cns_csa_n_shi0;
  output shr_mem_13_cns_csa_n_shi1;
  output shr_mem_13_cns_csb_n_shi0;
  output shr_mem_13_cns_csb_n_shi1;
  output [63:0] shr_mem_13_cns_dinb_shi0;
  output [63:0] shr_mem_13_cns_dinb_shi1;
  input [63:0] shr_mem_13_cns_douta_sho0;
  input [63:0] shr_mem_13_cns_douta_sho1;
  output shr_mem_13_cns_S1_pff;
  input din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_13_cns_S0_pff;


  // Interconnect Declarations
  reg dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_13_cns_PC0;
  reg shr_mem_13_cns_ppidx;
  reg [1:0] shr_mem_13_cns_ppown;
  wire shr_mem_13_cns_PC1;
  reg shr_mem_13_cns_ppidx_1;
  reg [1:0] shr_mem_13_cns_ppown_1;
  wire [6:0] shr_mem_13_shr_mem_13_mux_3_cse_pff;
  wire shr_mem_13_and_3_cse_pff;
  wire [1:0] shr_mem_13_acc_1_rmff;
  wire [3:0] nl_shr_mem_13_acc_1_rmff;
  wire shr_mem_13_xor_1_rmff;
  wire shr_mem_13_shr_mem_13_or_cse_pff;
  wire [1:0] shr_mem_13_acc_rmff;
  wire [3:0] nl_shr_mem_13_acc_rmff;
  wire shr_mem_13_xor_rmff;
  wire [6:0] shr_mem_13_shr_mem_13_mux_2_cse_pff;
  wire shr_mem_13_and_5_cse_pff;
  wire shr_mem_13_shr_mem_13_or_1_cse_pff;

  wire[0:0] shr_mem_13_mux_6_nl;
  wire[0:0] shr_mem_13_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_13_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_13_cns_R0;
  assign din_13_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_13_cns_R1;
  assign shr_mem_13_xor_rmff = shr_mem_13_cns_ppidx ^ shr_mem_13_cns_PC0;
  assign nl_shr_mem_13_acc_rmff = shr_mem_13_cns_ppown + conv_u2u_1_2(shr_mem_13_cns_PC0)
      + conv_s2u_1_2(shr_mem_13_cns_PC1);
  assign shr_mem_13_acc_rmff = nl_shr_mem_13_acc_rmff[1:0];
  assign shr_mem_13_cns_PC0 = shr_mem_13_cns_S0 & dout_13_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_13_xor_1_rmff = shr_mem_13_cns_ppidx_1 ^ shr_mem_13_cns_PC1;
  assign nl_shr_mem_13_acc_1_rmff = shr_mem_13_cns_ppown_1 + conv_u2u_1_2(shr_mem_13_cns_PC1)
      + conv_s2u_1_2(shr_mem_13_cns_PC0);
  assign shr_mem_13_acc_1_rmff = nl_shr_mem_13_acc_1_rmff[1:0];
  assign shr_mem_13_cns_PC1 = shr_mem_13_cns_S1 & din_13_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_13_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_13_cns_douta_sho0,
      shr_mem_13_cns_douta_sho1, shr_mem_13_cns_ppidx);
  assign din_13_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_13_cns_douta_sho0,
      shr_mem_13_cns_douta_sho1, shr_mem_13_cns_ppidx_1);
  assign shr_mem_13_cns_addra_shi0 = shr_mem_13_shr_mem_13_mux_3_cse_pff;
  assign shr_mem_13_cns_S1 = (shr_mem_13_cns_ppown_1!=2'b00);
  assign shr_mem_13_cns_S1_pff = (shr_mem_13_acc_1_rmff!=2'b00);
  assign shr_mem_13_and_3_cse_pff = shr_mem_13_cns_S1_pff & (~ shr_mem_13_xor_1_rmff);
  assign shr_mem_13_shr_mem_13_mux_3_cse_pff = MUX_v_7_2_2(dout_13_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_13_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_13_and_3_cse_pff);
  assign shr_mem_13_cns_addrb_shi0 = shr_mem_13_shr_mem_13_mux_3_cse_pff;
  assign shr_mem_13_cns_csa_n_shi0 = shr_mem_13_shr_mem_13_or_cse_pff;
  assign din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff =
      din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff =
      dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_13_cns_S0 = ~((shr_mem_13_cns_ppown==2'b10));
  assign shr_mem_13_cns_S0_pff = ~((shr_mem_13_acc_rmff==2'b10));
  assign shr_mem_13_mux_6_nl = MUX_s_1_2_2(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_13_and_3_cse_pff);
  assign shr_mem_13_shr_mem_13_or_cse_pff = (shr_mem_13_mux_6_nl) | (~((shr_mem_13_cns_S0_pff
      & (~ shr_mem_13_xor_rmff)) | shr_mem_13_and_3_cse_pff));
  assign shr_mem_13_cns_csb_n_shi0 = shr_mem_13_shr_mem_13_or_cse_pff;
  assign shr_mem_13_cns_dinb_shi0 = MUX_v_64_2_2(dout_13_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_13_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_13_and_3_cse_pff);
  assign shr_mem_13_cns_addra_shi1 = shr_mem_13_shr_mem_13_mux_2_cse_pff;
  assign shr_mem_13_and_5_cse_pff = shr_mem_13_cns_S1_pff & shr_mem_13_xor_1_rmff;
  assign shr_mem_13_shr_mem_13_mux_2_cse_pff = MUX_v_7_2_2(dout_13_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_13_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_13_and_5_cse_pff);
  assign shr_mem_13_cns_addrb_shi1 = shr_mem_13_shr_mem_13_mux_2_cse_pff;
  assign shr_mem_13_cns_csa_n_shi1 = shr_mem_13_shr_mem_13_or_1_cse_pff;
  assign shr_mem_13_mux_7_nl = MUX_s_1_2_2(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_13_and_5_cse_pff);
  assign shr_mem_13_shr_mem_13_or_1_cse_pff = (shr_mem_13_mux_7_nl) | (~((shr_mem_13_cns_S0_pff
      & shr_mem_13_xor_rmff) | shr_mem_13_and_5_cse_pff));
  assign shr_mem_13_cns_csb_n_shi1 = shr_mem_13_shr_mem_13_or_1_cse_pff;
  assign shr_mem_13_cns_dinb_shi1 = MUX_v_64_2_2(dout_13_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_13_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_13_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_13_cns_ppidx <= 1'b0;
      shr_mem_13_cns_ppown <= 2'b0;
      shr_mem_13_cns_ppidx_1 <= 1'b0;
      shr_mem_13_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_13_cns_ppidx <= shr_mem_13_xor_rmff;
      shr_mem_13_cns_ppown <= shr_mem_13_acc_rmff;
      shr_mem_13_cns_ppidx_1 <= shr_mem_13_xor_1_rmff;
      shr_mem_13_cns_ppown_1 <= shr_mem_13_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeoFsRV12_cns_bctl
// ------------------------------------------------------------------


module double_buffeoFsRV12_cns_bctl (
  clk, rst, dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_12_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_12_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_12_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_12_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_12_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_12_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_12_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_12_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_12_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_12_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_12_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_12_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_12_cns_S0, shr_mem_12_cns_R0, shr_mem_12_cns_S1, shr_mem_12_cns_R1,
      shr_mem_12_cns_addra_shi0, shr_mem_12_cns_addra_shi1, shr_mem_12_cns_addrb_shi0,
      shr_mem_12_cns_addrb_shi1, shr_mem_12_cns_csa_n_shi0, shr_mem_12_cns_csa_n_shi1,
      shr_mem_12_cns_csb_n_shi0, shr_mem_12_cns_csb_n_shi1, shr_mem_12_cns_dinb_shi0,
      shr_mem_12_cns_dinb_shi1, shr_mem_12_cns_douta_sho0, shr_mem_12_cns_douta_sho1,
      shr_mem_12_cns_S1_pff, din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_12_cns_S0_pff
);
  input clk;
  input rst;
  input dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_12_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_12_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_12_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_12_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_12_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_12_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_12_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_12_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_12_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_12_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_12_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_12_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_12_cns_S0;
  input shr_mem_12_cns_R0;
  output shr_mem_12_cns_S1;
  input shr_mem_12_cns_R1;
  output [6:0] shr_mem_12_cns_addra_shi0;
  output [6:0] shr_mem_12_cns_addra_shi1;
  output [6:0] shr_mem_12_cns_addrb_shi0;
  output [6:0] shr_mem_12_cns_addrb_shi1;
  output shr_mem_12_cns_csa_n_shi0;
  output shr_mem_12_cns_csa_n_shi1;
  output shr_mem_12_cns_csb_n_shi0;
  output shr_mem_12_cns_csb_n_shi1;
  output [63:0] shr_mem_12_cns_dinb_shi0;
  output [63:0] shr_mem_12_cns_dinb_shi1;
  input [63:0] shr_mem_12_cns_douta_sho0;
  input [63:0] shr_mem_12_cns_douta_sho1;
  output shr_mem_12_cns_S1_pff;
  input din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_12_cns_S0_pff;


  // Interconnect Declarations
  reg dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_12_cns_PC0;
  reg shr_mem_12_cns_ppidx;
  reg [1:0] shr_mem_12_cns_ppown;
  wire shr_mem_12_cns_PC1;
  reg shr_mem_12_cns_ppidx_1;
  reg [1:0] shr_mem_12_cns_ppown_1;
  wire [6:0] shr_mem_12_shr_mem_12_mux_3_cse_pff;
  wire shr_mem_12_and_3_cse_pff;
  wire [1:0] shr_mem_12_acc_1_rmff;
  wire [3:0] nl_shr_mem_12_acc_1_rmff;
  wire shr_mem_12_xor_1_rmff;
  wire shr_mem_12_shr_mem_12_or_cse_pff;
  wire [1:0] shr_mem_12_acc_rmff;
  wire [3:0] nl_shr_mem_12_acc_rmff;
  wire shr_mem_12_xor_rmff;
  wire [6:0] shr_mem_12_shr_mem_12_mux_2_cse_pff;
  wire shr_mem_12_and_5_cse_pff;
  wire shr_mem_12_shr_mem_12_or_1_cse_pff;

  wire[0:0] shr_mem_12_mux_6_nl;
  wire[0:0] shr_mem_12_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_12_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_12_cns_R0;
  assign din_12_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_12_cns_R1;
  assign shr_mem_12_xor_rmff = shr_mem_12_cns_ppidx ^ shr_mem_12_cns_PC0;
  assign nl_shr_mem_12_acc_rmff = shr_mem_12_cns_ppown + conv_u2u_1_2(shr_mem_12_cns_PC0)
      + conv_s2u_1_2(shr_mem_12_cns_PC1);
  assign shr_mem_12_acc_rmff = nl_shr_mem_12_acc_rmff[1:0];
  assign shr_mem_12_cns_PC0 = shr_mem_12_cns_S0 & dout_12_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_12_xor_1_rmff = shr_mem_12_cns_ppidx_1 ^ shr_mem_12_cns_PC1;
  assign nl_shr_mem_12_acc_1_rmff = shr_mem_12_cns_ppown_1 + conv_u2u_1_2(shr_mem_12_cns_PC1)
      + conv_s2u_1_2(shr_mem_12_cns_PC0);
  assign shr_mem_12_acc_1_rmff = nl_shr_mem_12_acc_1_rmff[1:0];
  assign shr_mem_12_cns_PC1 = shr_mem_12_cns_S1 & din_12_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_12_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_12_cns_douta_sho0,
      shr_mem_12_cns_douta_sho1, shr_mem_12_cns_ppidx);
  assign din_12_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_12_cns_douta_sho0,
      shr_mem_12_cns_douta_sho1, shr_mem_12_cns_ppidx_1);
  assign shr_mem_12_cns_addra_shi0 = shr_mem_12_shr_mem_12_mux_3_cse_pff;
  assign shr_mem_12_cns_S1 = (shr_mem_12_cns_ppown_1!=2'b00);
  assign shr_mem_12_cns_S1_pff = (shr_mem_12_acc_1_rmff!=2'b00);
  assign shr_mem_12_and_3_cse_pff = shr_mem_12_cns_S1_pff & (~ shr_mem_12_xor_1_rmff);
  assign shr_mem_12_shr_mem_12_mux_3_cse_pff = MUX_v_7_2_2(dout_12_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_12_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_12_and_3_cse_pff);
  assign shr_mem_12_cns_addrb_shi0 = shr_mem_12_shr_mem_12_mux_3_cse_pff;
  assign shr_mem_12_cns_csa_n_shi0 = shr_mem_12_shr_mem_12_or_cse_pff;
  assign din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff =
      din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff =
      dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_12_cns_S0 = ~((shr_mem_12_cns_ppown==2'b10));
  assign shr_mem_12_cns_S0_pff = ~((shr_mem_12_acc_rmff==2'b10));
  assign shr_mem_12_mux_6_nl = MUX_s_1_2_2(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_12_and_3_cse_pff);
  assign shr_mem_12_shr_mem_12_or_cse_pff = (shr_mem_12_mux_6_nl) | (~((shr_mem_12_cns_S0_pff
      & (~ shr_mem_12_xor_rmff)) | shr_mem_12_and_3_cse_pff));
  assign shr_mem_12_cns_csb_n_shi0 = shr_mem_12_shr_mem_12_or_cse_pff;
  assign shr_mem_12_cns_dinb_shi0 = MUX_v_64_2_2(dout_12_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_12_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_12_and_3_cse_pff);
  assign shr_mem_12_cns_addra_shi1 = shr_mem_12_shr_mem_12_mux_2_cse_pff;
  assign shr_mem_12_and_5_cse_pff = shr_mem_12_cns_S1_pff & shr_mem_12_xor_1_rmff;
  assign shr_mem_12_shr_mem_12_mux_2_cse_pff = MUX_v_7_2_2(dout_12_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_12_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_12_and_5_cse_pff);
  assign shr_mem_12_cns_addrb_shi1 = shr_mem_12_shr_mem_12_mux_2_cse_pff;
  assign shr_mem_12_cns_csa_n_shi1 = shr_mem_12_shr_mem_12_or_1_cse_pff;
  assign shr_mem_12_mux_7_nl = MUX_s_1_2_2(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_12_and_5_cse_pff);
  assign shr_mem_12_shr_mem_12_or_1_cse_pff = (shr_mem_12_mux_7_nl) | (~((shr_mem_12_cns_S0_pff
      & shr_mem_12_xor_rmff) | shr_mem_12_and_5_cse_pff));
  assign shr_mem_12_cns_csb_n_shi1 = shr_mem_12_shr_mem_12_or_1_cse_pff;
  assign shr_mem_12_cns_dinb_shi1 = MUX_v_64_2_2(dout_12_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_12_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_12_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_12_cns_ppidx <= 1'b0;
      shr_mem_12_cns_ppown <= 2'b0;
      shr_mem_12_cns_ppidx_1 <= 1'b0;
      shr_mem_12_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_12_cns_ppidx <= shr_mem_12_xor_rmff;
      shr_mem_12_cns_ppown <= shr_mem_12_acc_rmff;
      shr_mem_12_cns_ppidx_1 <= shr_mem_12_xor_1_rmff;
      shr_mem_12_cns_ppown_1 <= shr_mem_12_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeoFsRV11_cns_bctl
// ------------------------------------------------------------------


module double_buffeoFsRV11_cns_bctl (
  clk, rst, dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_11_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_11_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_11_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_11_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_11_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_11_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_11_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_11_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_11_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_11_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_11_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_11_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_11_cns_S0, shr_mem_11_cns_R0, shr_mem_11_cns_S1, shr_mem_11_cns_R1,
      shr_mem_11_cns_addra_shi0, shr_mem_11_cns_addra_shi1, shr_mem_11_cns_addrb_shi0,
      shr_mem_11_cns_addrb_shi1, shr_mem_11_cns_csa_n_shi0, shr_mem_11_cns_csa_n_shi1,
      shr_mem_11_cns_csb_n_shi0, shr_mem_11_cns_csb_n_shi1, shr_mem_11_cns_dinb_shi0,
      shr_mem_11_cns_dinb_shi1, shr_mem_11_cns_douta_sho0, shr_mem_11_cns_douta_sho1,
      shr_mem_11_cns_S1_pff, din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_11_cns_S0_pff
);
  input clk;
  input rst;
  input dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_11_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_11_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_11_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_11_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_11_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_11_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_11_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_11_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_11_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_11_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_11_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_11_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_11_cns_S0;
  input shr_mem_11_cns_R0;
  output shr_mem_11_cns_S1;
  input shr_mem_11_cns_R1;
  output [6:0] shr_mem_11_cns_addra_shi0;
  output [6:0] shr_mem_11_cns_addra_shi1;
  output [6:0] shr_mem_11_cns_addrb_shi0;
  output [6:0] shr_mem_11_cns_addrb_shi1;
  output shr_mem_11_cns_csa_n_shi0;
  output shr_mem_11_cns_csa_n_shi1;
  output shr_mem_11_cns_csb_n_shi0;
  output shr_mem_11_cns_csb_n_shi1;
  output [63:0] shr_mem_11_cns_dinb_shi0;
  output [63:0] shr_mem_11_cns_dinb_shi1;
  input [63:0] shr_mem_11_cns_douta_sho0;
  input [63:0] shr_mem_11_cns_douta_sho1;
  output shr_mem_11_cns_S1_pff;
  input din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_11_cns_S0_pff;


  // Interconnect Declarations
  reg dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_11_cns_PC0;
  reg shr_mem_11_cns_ppidx;
  reg [1:0] shr_mem_11_cns_ppown;
  wire shr_mem_11_cns_PC1;
  reg shr_mem_11_cns_ppidx_1;
  reg [1:0] shr_mem_11_cns_ppown_1;
  wire [6:0] shr_mem_11_shr_mem_11_mux_3_cse_pff;
  wire shr_mem_11_and_3_cse_pff;
  wire [1:0] shr_mem_11_acc_1_rmff;
  wire [3:0] nl_shr_mem_11_acc_1_rmff;
  wire shr_mem_11_xor_1_rmff;
  wire shr_mem_11_shr_mem_11_or_cse_pff;
  wire [1:0] shr_mem_11_acc_rmff;
  wire [3:0] nl_shr_mem_11_acc_rmff;
  wire shr_mem_11_xor_rmff;
  wire [6:0] shr_mem_11_shr_mem_11_mux_2_cse_pff;
  wire shr_mem_11_and_5_cse_pff;
  wire shr_mem_11_shr_mem_11_or_1_cse_pff;

  wire[0:0] shr_mem_11_mux_6_nl;
  wire[0:0] shr_mem_11_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_11_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_11_cns_R0;
  assign din_11_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_11_cns_R1;
  assign shr_mem_11_xor_rmff = shr_mem_11_cns_ppidx ^ shr_mem_11_cns_PC0;
  assign nl_shr_mem_11_acc_rmff = shr_mem_11_cns_ppown + conv_u2u_1_2(shr_mem_11_cns_PC0)
      + conv_s2u_1_2(shr_mem_11_cns_PC1);
  assign shr_mem_11_acc_rmff = nl_shr_mem_11_acc_rmff[1:0];
  assign shr_mem_11_cns_PC0 = shr_mem_11_cns_S0 & dout_11_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_11_xor_1_rmff = shr_mem_11_cns_ppidx_1 ^ shr_mem_11_cns_PC1;
  assign nl_shr_mem_11_acc_1_rmff = shr_mem_11_cns_ppown_1 + conv_u2u_1_2(shr_mem_11_cns_PC1)
      + conv_s2u_1_2(shr_mem_11_cns_PC0);
  assign shr_mem_11_acc_1_rmff = nl_shr_mem_11_acc_1_rmff[1:0];
  assign shr_mem_11_cns_PC1 = shr_mem_11_cns_S1 & din_11_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_11_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_11_cns_douta_sho0,
      shr_mem_11_cns_douta_sho1, shr_mem_11_cns_ppidx);
  assign din_11_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_11_cns_douta_sho0,
      shr_mem_11_cns_douta_sho1, shr_mem_11_cns_ppidx_1);
  assign shr_mem_11_cns_addra_shi0 = shr_mem_11_shr_mem_11_mux_3_cse_pff;
  assign shr_mem_11_cns_S1 = (shr_mem_11_cns_ppown_1!=2'b00);
  assign shr_mem_11_cns_S1_pff = (shr_mem_11_acc_1_rmff!=2'b00);
  assign shr_mem_11_and_3_cse_pff = shr_mem_11_cns_S1_pff & (~ shr_mem_11_xor_1_rmff);
  assign shr_mem_11_shr_mem_11_mux_3_cse_pff = MUX_v_7_2_2(dout_11_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_11_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_11_and_3_cse_pff);
  assign shr_mem_11_cns_addrb_shi0 = shr_mem_11_shr_mem_11_mux_3_cse_pff;
  assign shr_mem_11_cns_csa_n_shi0 = shr_mem_11_shr_mem_11_or_cse_pff;
  assign din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff =
      din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff =
      dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_11_cns_S0 = ~((shr_mem_11_cns_ppown==2'b10));
  assign shr_mem_11_cns_S0_pff = ~((shr_mem_11_acc_rmff==2'b10));
  assign shr_mem_11_mux_6_nl = MUX_s_1_2_2(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_11_and_3_cse_pff);
  assign shr_mem_11_shr_mem_11_or_cse_pff = (shr_mem_11_mux_6_nl) | (~((shr_mem_11_cns_S0_pff
      & (~ shr_mem_11_xor_rmff)) | shr_mem_11_and_3_cse_pff));
  assign shr_mem_11_cns_csb_n_shi0 = shr_mem_11_shr_mem_11_or_cse_pff;
  assign shr_mem_11_cns_dinb_shi0 = MUX_v_64_2_2(dout_11_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_11_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_11_and_3_cse_pff);
  assign shr_mem_11_cns_addra_shi1 = shr_mem_11_shr_mem_11_mux_2_cse_pff;
  assign shr_mem_11_and_5_cse_pff = shr_mem_11_cns_S1_pff & shr_mem_11_xor_1_rmff;
  assign shr_mem_11_shr_mem_11_mux_2_cse_pff = MUX_v_7_2_2(dout_11_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_11_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_11_and_5_cse_pff);
  assign shr_mem_11_cns_addrb_shi1 = shr_mem_11_shr_mem_11_mux_2_cse_pff;
  assign shr_mem_11_cns_csa_n_shi1 = shr_mem_11_shr_mem_11_or_1_cse_pff;
  assign shr_mem_11_mux_7_nl = MUX_s_1_2_2(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_11_and_5_cse_pff);
  assign shr_mem_11_shr_mem_11_or_1_cse_pff = (shr_mem_11_mux_7_nl) | (~((shr_mem_11_cns_S0_pff
      & shr_mem_11_xor_rmff) | shr_mem_11_and_5_cse_pff));
  assign shr_mem_11_cns_csb_n_shi1 = shr_mem_11_shr_mem_11_or_1_cse_pff;
  assign shr_mem_11_cns_dinb_shi1 = MUX_v_64_2_2(dout_11_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_11_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_11_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_11_cns_ppidx <= 1'b0;
      shr_mem_11_cns_ppown <= 2'b0;
      shr_mem_11_cns_ppidx_1 <= 1'b0;
      shr_mem_11_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_11_cns_ppidx <= shr_mem_11_xor_rmff;
      shr_mem_11_cns_ppown <= shr_mem_11_acc_rmff;
      shr_mem_11_cns_ppidx_1 <= shr_mem_11_xor_1_rmff;
      shr_mem_11_cns_ppown_1 <= shr_mem_11_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeoFsRV10_cns_bctl
// ------------------------------------------------------------------


module double_buffeoFsRV10_cns_bctl (
  clk, rst, dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_10_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_10_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_10_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_10_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_10_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_10_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_10_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_10_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_10_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_10_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_10_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_10_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_10_cns_S0, shr_mem_10_cns_R0, shr_mem_10_cns_S1, shr_mem_10_cns_R1,
      shr_mem_10_cns_addra_shi0, shr_mem_10_cns_addra_shi1, shr_mem_10_cns_addrb_shi0,
      shr_mem_10_cns_addrb_shi1, shr_mem_10_cns_csa_n_shi0, shr_mem_10_cns_csa_n_shi1,
      shr_mem_10_cns_csb_n_shi0, shr_mem_10_cns_csb_n_shi1, shr_mem_10_cns_dinb_shi0,
      shr_mem_10_cns_dinb_shi1, shr_mem_10_cns_douta_sho0, shr_mem_10_cns_douta_sho1,
      shr_mem_10_cns_S1_pff, din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_10_cns_S0_pff
);
  input clk;
  input rst;
  input dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_10_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_10_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_10_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_10_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_10_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_10_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_10_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_10_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_10_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_10_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_10_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_10_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_10_cns_S0;
  input shr_mem_10_cns_R0;
  output shr_mem_10_cns_S1;
  input shr_mem_10_cns_R1;
  output [6:0] shr_mem_10_cns_addra_shi0;
  output [6:0] shr_mem_10_cns_addra_shi1;
  output [6:0] shr_mem_10_cns_addrb_shi0;
  output [6:0] shr_mem_10_cns_addrb_shi1;
  output shr_mem_10_cns_csa_n_shi0;
  output shr_mem_10_cns_csa_n_shi1;
  output shr_mem_10_cns_csb_n_shi0;
  output shr_mem_10_cns_csb_n_shi1;
  output [63:0] shr_mem_10_cns_dinb_shi0;
  output [63:0] shr_mem_10_cns_dinb_shi1;
  input [63:0] shr_mem_10_cns_douta_sho0;
  input [63:0] shr_mem_10_cns_douta_sho1;
  output shr_mem_10_cns_S1_pff;
  input din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_10_cns_S0_pff;


  // Interconnect Declarations
  reg dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_10_cns_PC0;
  reg shr_mem_10_cns_ppidx;
  reg [1:0] shr_mem_10_cns_ppown;
  wire shr_mem_10_cns_PC1;
  reg shr_mem_10_cns_ppidx_1;
  reg [1:0] shr_mem_10_cns_ppown_1;
  wire [6:0] shr_mem_10_shr_mem_10_mux_3_cse_pff;
  wire shr_mem_10_and_3_cse_pff;
  wire [1:0] shr_mem_10_acc_1_rmff;
  wire [3:0] nl_shr_mem_10_acc_1_rmff;
  wire shr_mem_10_xor_1_rmff;
  wire shr_mem_10_shr_mem_10_or_cse_pff;
  wire [1:0] shr_mem_10_acc_rmff;
  wire [3:0] nl_shr_mem_10_acc_rmff;
  wire shr_mem_10_xor_rmff;
  wire [6:0] shr_mem_10_shr_mem_10_mux_2_cse_pff;
  wire shr_mem_10_and_5_cse_pff;
  wire shr_mem_10_shr_mem_10_or_1_cse_pff;

  wire[0:0] shr_mem_10_mux_6_nl;
  wire[0:0] shr_mem_10_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_10_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_10_cns_R0;
  assign din_10_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_10_cns_R1;
  assign shr_mem_10_xor_rmff = shr_mem_10_cns_ppidx ^ shr_mem_10_cns_PC0;
  assign nl_shr_mem_10_acc_rmff = shr_mem_10_cns_ppown + conv_u2u_1_2(shr_mem_10_cns_PC0)
      + conv_s2u_1_2(shr_mem_10_cns_PC1);
  assign shr_mem_10_acc_rmff = nl_shr_mem_10_acc_rmff[1:0];
  assign shr_mem_10_cns_PC0 = shr_mem_10_cns_S0 & dout_10_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_10_xor_1_rmff = shr_mem_10_cns_ppidx_1 ^ shr_mem_10_cns_PC1;
  assign nl_shr_mem_10_acc_1_rmff = shr_mem_10_cns_ppown_1 + conv_u2u_1_2(shr_mem_10_cns_PC1)
      + conv_s2u_1_2(shr_mem_10_cns_PC0);
  assign shr_mem_10_acc_1_rmff = nl_shr_mem_10_acc_1_rmff[1:0];
  assign shr_mem_10_cns_PC1 = shr_mem_10_cns_S1 & din_10_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_10_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_10_cns_douta_sho0,
      shr_mem_10_cns_douta_sho1, shr_mem_10_cns_ppidx);
  assign din_10_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_10_cns_douta_sho0,
      shr_mem_10_cns_douta_sho1, shr_mem_10_cns_ppidx_1);
  assign shr_mem_10_cns_addra_shi0 = shr_mem_10_shr_mem_10_mux_3_cse_pff;
  assign shr_mem_10_cns_S1 = (shr_mem_10_cns_ppown_1!=2'b00);
  assign shr_mem_10_cns_S1_pff = (shr_mem_10_acc_1_rmff!=2'b00);
  assign shr_mem_10_and_3_cse_pff = shr_mem_10_cns_S1_pff & (~ shr_mem_10_xor_1_rmff);
  assign shr_mem_10_shr_mem_10_mux_3_cse_pff = MUX_v_7_2_2(dout_10_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_10_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_10_and_3_cse_pff);
  assign shr_mem_10_cns_addrb_shi0 = shr_mem_10_shr_mem_10_mux_3_cse_pff;
  assign shr_mem_10_cns_csa_n_shi0 = shr_mem_10_shr_mem_10_or_cse_pff;
  assign din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff =
      din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff =
      dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_10_cns_S0 = ~((shr_mem_10_cns_ppown==2'b10));
  assign shr_mem_10_cns_S0_pff = ~((shr_mem_10_acc_rmff==2'b10));
  assign shr_mem_10_mux_6_nl = MUX_s_1_2_2(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_10_and_3_cse_pff);
  assign shr_mem_10_shr_mem_10_or_cse_pff = (shr_mem_10_mux_6_nl) | (~((shr_mem_10_cns_S0_pff
      & (~ shr_mem_10_xor_rmff)) | shr_mem_10_and_3_cse_pff));
  assign shr_mem_10_cns_csb_n_shi0 = shr_mem_10_shr_mem_10_or_cse_pff;
  assign shr_mem_10_cns_dinb_shi0 = MUX_v_64_2_2(dout_10_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_10_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_10_and_3_cse_pff);
  assign shr_mem_10_cns_addra_shi1 = shr_mem_10_shr_mem_10_mux_2_cse_pff;
  assign shr_mem_10_and_5_cse_pff = shr_mem_10_cns_S1_pff & shr_mem_10_xor_1_rmff;
  assign shr_mem_10_shr_mem_10_mux_2_cse_pff = MUX_v_7_2_2(dout_10_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_10_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_10_and_5_cse_pff);
  assign shr_mem_10_cns_addrb_shi1 = shr_mem_10_shr_mem_10_mux_2_cse_pff;
  assign shr_mem_10_cns_csa_n_shi1 = shr_mem_10_shr_mem_10_or_1_cse_pff;
  assign shr_mem_10_mux_7_nl = MUX_s_1_2_2(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_10_and_5_cse_pff);
  assign shr_mem_10_shr_mem_10_or_1_cse_pff = (shr_mem_10_mux_7_nl) | (~((shr_mem_10_cns_S0_pff
      & shr_mem_10_xor_rmff) | shr_mem_10_and_5_cse_pff));
  assign shr_mem_10_cns_csb_n_shi1 = shr_mem_10_shr_mem_10_or_1_cse_pff;
  assign shr_mem_10_cns_dinb_shi1 = MUX_v_64_2_2(dout_10_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_10_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_10_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_10_cns_ppidx <= 1'b0;
      shr_mem_10_cns_ppown <= 2'b0;
      shr_mem_10_cns_ppidx_1 <= 1'b0;
      shr_mem_10_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_10_cns_ppidx <= shr_mem_10_xor_rmff;
      shr_mem_10_cns_ppown <= shr_mem_10_acc_rmff;
      shr_mem_10_cns_ppidx_1 <= shr_mem_10_xor_1_rmff;
      shr_mem_10_cns_ppown_1 <= shr_mem_10_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeaIgYu_9_cns_bctl
// ------------------------------------------------------------------


module double_buffeaIgYu_9_cns_bctl (
  clk, rst, dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_9_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_9_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_9_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_9_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_9_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_9_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_9_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_9_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_9_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_9_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_9_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_9_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_9_cns_S0, shr_mem_9_cns_R0, shr_mem_9_cns_S1, shr_mem_9_cns_R1, shr_mem_9_cns_addra_shi0,
      shr_mem_9_cns_addra_shi1, shr_mem_9_cns_addrb_shi0, shr_mem_9_cns_addrb_shi1,
      shr_mem_9_cns_csa_n_shi0, shr_mem_9_cns_csa_n_shi1, shr_mem_9_cns_csb_n_shi0,
      shr_mem_9_cns_csb_n_shi1, shr_mem_9_cns_dinb_shi0, shr_mem_9_cns_dinb_shi1,
      shr_mem_9_cns_douta_sho0, shr_mem_9_cns_douta_sho1, shr_mem_9_cns_S1_pff, din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_9_cns_S0_pff
);
  input clk;
  input rst;
  input dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_9_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_9_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_9_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_9_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_9_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_9_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_9_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_9_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_9_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_9_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_9_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_9_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_9_cns_S0;
  input shr_mem_9_cns_R0;
  output shr_mem_9_cns_S1;
  input shr_mem_9_cns_R1;
  output [6:0] shr_mem_9_cns_addra_shi0;
  output [6:0] shr_mem_9_cns_addra_shi1;
  output [6:0] shr_mem_9_cns_addrb_shi0;
  output [6:0] shr_mem_9_cns_addrb_shi1;
  output shr_mem_9_cns_csa_n_shi0;
  output shr_mem_9_cns_csa_n_shi1;
  output shr_mem_9_cns_csb_n_shi0;
  output shr_mem_9_cns_csb_n_shi1;
  output [63:0] shr_mem_9_cns_dinb_shi0;
  output [63:0] shr_mem_9_cns_dinb_shi1;
  input [63:0] shr_mem_9_cns_douta_sho0;
  input [63:0] shr_mem_9_cns_douta_sho1;
  output shr_mem_9_cns_S1_pff;
  input din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_9_cns_S0_pff;


  // Interconnect Declarations
  reg dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_9_cns_PC0;
  reg shr_mem_9_cns_ppidx;
  reg [1:0] shr_mem_9_cns_ppown;
  wire shr_mem_9_cns_PC1;
  reg shr_mem_9_cns_ppidx_1;
  reg [1:0] shr_mem_9_cns_ppown_1;
  wire [6:0] shr_mem_9_shr_mem_9_mux_3_cse_pff;
  wire shr_mem_9_and_3_cse_pff;
  wire [1:0] shr_mem_9_acc_1_rmff;
  wire [3:0] nl_shr_mem_9_acc_1_rmff;
  wire shr_mem_9_xor_1_rmff;
  wire shr_mem_9_shr_mem_9_or_cse_pff;
  wire [1:0] shr_mem_9_acc_rmff;
  wire [3:0] nl_shr_mem_9_acc_rmff;
  wire shr_mem_9_xor_rmff;
  wire [6:0] shr_mem_9_shr_mem_9_mux_2_cse_pff;
  wire shr_mem_9_and_5_cse_pff;
  wire shr_mem_9_shr_mem_9_or_1_cse_pff;

  wire[0:0] shr_mem_9_mux_6_nl;
  wire[0:0] shr_mem_9_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_9_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_9_cns_R0;
  assign din_9_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_9_cns_R1;
  assign shr_mem_9_xor_rmff = shr_mem_9_cns_ppidx ^ shr_mem_9_cns_PC0;
  assign nl_shr_mem_9_acc_rmff = shr_mem_9_cns_ppown + conv_u2u_1_2(shr_mem_9_cns_PC0)
      + conv_s2u_1_2(shr_mem_9_cns_PC1);
  assign shr_mem_9_acc_rmff = nl_shr_mem_9_acc_rmff[1:0];
  assign shr_mem_9_cns_PC0 = shr_mem_9_cns_S0 & dout_9_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_9_xor_1_rmff = shr_mem_9_cns_ppidx_1 ^ shr_mem_9_cns_PC1;
  assign nl_shr_mem_9_acc_1_rmff = shr_mem_9_cns_ppown_1 + conv_u2u_1_2(shr_mem_9_cns_PC1)
      + conv_s2u_1_2(shr_mem_9_cns_PC0);
  assign shr_mem_9_acc_1_rmff = nl_shr_mem_9_acc_1_rmff[1:0];
  assign shr_mem_9_cns_PC1 = shr_mem_9_cns_S1 & din_9_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_9_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_9_cns_douta_sho0,
      shr_mem_9_cns_douta_sho1, shr_mem_9_cns_ppidx);
  assign din_9_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_9_cns_douta_sho0,
      shr_mem_9_cns_douta_sho1, shr_mem_9_cns_ppidx_1);
  assign shr_mem_9_cns_addra_shi0 = shr_mem_9_shr_mem_9_mux_3_cse_pff;
  assign shr_mem_9_cns_S1 = (shr_mem_9_cns_ppown_1!=2'b00);
  assign shr_mem_9_cns_S1_pff = (shr_mem_9_acc_1_rmff!=2'b00);
  assign shr_mem_9_and_3_cse_pff = shr_mem_9_cns_S1_pff & (~ shr_mem_9_xor_1_rmff);
  assign shr_mem_9_shr_mem_9_mux_3_cse_pff = MUX_v_7_2_2(dout_9_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_9_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_9_and_3_cse_pff);
  assign shr_mem_9_cns_addrb_shi0 = shr_mem_9_shr_mem_9_mux_3_cse_pff;
  assign shr_mem_9_cns_csa_n_shi0 = shr_mem_9_shr_mem_9_or_cse_pff;
  assign din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff = din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff = dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_9_cns_S0 = ~((shr_mem_9_cns_ppown==2'b10));
  assign shr_mem_9_cns_S0_pff = ~((shr_mem_9_acc_rmff==2'b10));
  assign shr_mem_9_mux_6_nl = MUX_s_1_2_2(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_9_and_3_cse_pff);
  assign shr_mem_9_shr_mem_9_or_cse_pff = (shr_mem_9_mux_6_nl) | (~((shr_mem_9_cns_S0_pff
      & (~ shr_mem_9_xor_rmff)) | shr_mem_9_and_3_cse_pff));
  assign shr_mem_9_cns_csb_n_shi0 = shr_mem_9_shr_mem_9_or_cse_pff;
  assign shr_mem_9_cns_dinb_shi0 = MUX_v_64_2_2(dout_9_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_9_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_9_and_3_cse_pff);
  assign shr_mem_9_cns_addra_shi1 = shr_mem_9_shr_mem_9_mux_2_cse_pff;
  assign shr_mem_9_and_5_cse_pff = shr_mem_9_cns_S1_pff & shr_mem_9_xor_1_rmff;
  assign shr_mem_9_shr_mem_9_mux_2_cse_pff = MUX_v_7_2_2(dout_9_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_9_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_9_and_5_cse_pff);
  assign shr_mem_9_cns_addrb_shi1 = shr_mem_9_shr_mem_9_mux_2_cse_pff;
  assign shr_mem_9_cns_csa_n_shi1 = shr_mem_9_shr_mem_9_or_1_cse_pff;
  assign shr_mem_9_mux_7_nl = MUX_s_1_2_2(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_9_and_5_cse_pff);
  assign shr_mem_9_shr_mem_9_or_1_cse_pff = (shr_mem_9_mux_7_nl) | (~((shr_mem_9_cns_S0_pff
      & shr_mem_9_xor_rmff) | shr_mem_9_and_5_cse_pff));
  assign shr_mem_9_cns_csb_n_shi1 = shr_mem_9_shr_mem_9_or_1_cse_pff;
  assign shr_mem_9_cns_dinb_shi1 = MUX_v_64_2_2(dout_9_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_9_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_9_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_9_cns_ppidx <= 1'b0;
      shr_mem_9_cns_ppown <= 2'b0;
      shr_mem_9_cns_ppidx_1 <= 1'b0;
      shr_mem_9_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_9_cns_ppidx <= shr_mem_9_xor_rmff;
      shr_mem_9_cns_ppown <= shr_mem_9_acc_rmff;
      shr_mem_9_cns_ppidx_1 <= shr_mem_9_xor_1_rmff;
      shr_mem_9_cns_ppown_1 <= shr_mem_9_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeaIgYu_8_cns_bctl
// ------------------------------------------------------------------


module double_buffeaIgYu_8_cns_bctl (
  clk, rst, dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_8_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_8_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_8_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_8_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_8_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_8_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_8_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_8_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_8_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_8_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_8_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_8_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_8_cns_S0, shr_mem_8_cns_R0, shr_mem_8_cns_S1, shr_mem_8_cns_R1, shr_mem_8_cns_addra_shi0,
      shr_mem_8_cns_addra_shi1, shr_mem_8_cns_addrb_shi0, shr_mem_8_cns_addrb_shi1,
      shr_mem_8_cns_csa_n_shi0, shr_mem_8_cns_csa_n_shi1, shr_mem_8_cns_csb_n_shi0,
      shr_mem_8_cns_csb_n_shi1, shr_mem_8_cns_dinb_shi0, shr_mem_8_cns_dinb_shi1,
      shr_mem_8_cns_douta_sho0, shr_mem_8_cns_douta_sho1, shr_mem_8_cns_S1_pff, din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_8_cns_S0_pff
);
  input clk;
  input rst;
  input dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_8_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_8_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_8_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_8_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_8_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_8_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_8_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_8_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_8_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_8_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_8_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_8_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_8_cns_S0;
  input shr_mem_8_cns_R0;
  output shr_mem_8_cns_S1;
  input shr_mem_8_cns_R1;
  output [6:0] shr_mem_8_cns_addra_shi0;
  output [6:0] shr_mem_8_cns_addra_shi1;
  output [6:0] shr_mem_8_cns_addrb_shi0;
  output [6:0] shr_mem_8_cns_addrb_shi1;
  output shr_mem_8_cns_csa_n_shi0;
  output shr_mem_8_cns_csa_n_shi1;
  output shr_mem_8_cns_csb_n_shi0;
  output shr_mem_8_cns_csb_n_shi1;
  output [63:0] shr_mem_8_cns_dinb_shi0;
  output [63:0] shr_mem_8_cns_dinb_shi1;
  input [63:0] shr_mem_8_cns_douta_sho0;
  input [63:0] shr_mem_8_cns_douta_sho1;
  output shr_mem_8_cns_S1_pff;
  input din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_8_cns_S0_pff;


  // Interconnect Declarations
  reg dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_8_cns_PC0;
  reg shr_mem_8_cns_ppidx;
  reg [1:0] shr_mem_8_cns_ppown;
  wire shr_mem_8_cns_PC1;
  reg shr_mem_8_cns_ppidx_1;
  reg [1:0] shr_mem_8_cns_ppown_1;
  wire [6:0] shr_mem_8_shr_mem_8_mux_3_cse_pff;
  wire shr_mem_8_and_3_cse_pff;
  wire [1:0] shr_mem_8_acc_1_rmff;
  wire [3:0] nl_shr_mem_8_acc_1_rmff;
  wire shr_mem_8_xor_1_rmff;
  wire shr_mem_8_shr_mem_8_or_cse_pff;
  wire [1:0] shr_mem_8_acc_rmff;
  wire [3:0] nl_shr_mem_8_acc_rmff;
  wire shr_mem_8_xor_rmff;
  wire [6:0] shr_mem_8_shr_mem_8_mux_2_cse_pff;
  wire shr_mem_8_and_5_cse_pff;
  wire shr_mem_8_shr_mem_8_or_1_cse_pff;

  wire[0:0] shr_mem_8_mux_6_nl;
  wire[0:0] shr_mem_8_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_8_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_8_cns_R0;
  assign din_8_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_8_cns_R1;
  assign shr_mem_8_xor_rmff = shr_mem_8_cns_ppidx ^ shr_mem_8_cns_PC0;
  assign nl_shr_mem_8_acc_rmff = shr_mem_8_cns_ppown + conv_u2u_1_2(shr_mem_8_cns_PC0)
      + conv_s2u_1_2(shr_mem_8_cns_PC1);
  assign shr_mem_8_acc_rmff = nl_shr_mem_8_acc_rmff[1:0];
  assign shr_mem_8_cns_PC0 = shr_mem_8_cns_S0 & dout_8_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_8_xor_1_rmff = shr_mem_8_cns_ppidx_1 ^ shr_mem_8_cns_PC1;
  assign nl_shr_mem_8_acc_1_rmff = shr_mem_8_cns_ppown_1 + conv_u2u_1_2(shr_mem_8_cns_PC1)
      + conv_s2u_1_2(shr_mem_8_cns_PC0);
  assign shr_mem_8_acc_1_rmff = nl_shr_mem_8_acc_1_rmff[1:0];
  assign shr_mem_8_cns_PC1 = shr_mem_8_cns_S1 & din_8_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_8_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_8_cns_douta_sho0,
      shr_mem_8_cns_douta_sho1, shr_mem_8_cns_ppidx);
  assign din_8_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_8_cns_douta_sho0,
      shr_mem_8_cns_douta_sho1, shr_mem_8_cns_ppidx_1);
  assign shr_mem_8_cns_addra_shi0 = shr_mem_8_shr_mem_8_mux_3_cse_pff;
  assign shr_mem_8_cns_S1 = (shr_mem_8_cns_ppown_1!=2'b00);
  assign shr_mem_8_cns_S1_pff = (shr_mem_8_acc_1_rmff!=2'b00);
  assign shr_mem_8_and_3_cse_pff = shr_mem_8_cns_S1_pff & (~ shr_mem_8_xor_1_rmff);
  assign shr_mem_8_shr_mem_8_mux_3_cse_pff = MUX_v_7_2_2(dout_8_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_8_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_8_and_3_cse_pff);
  assign shr_mem_8_cns_addrb_shi0 = shr_mem_8_shr_mem_8_mux_3_cse_pff;
  assign shr_mem_8_cns_csa_n_shi0 = shr_mem_8_shr_mem_8_or_cse_pff;
  assign din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff = din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff = dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_8_cns_S0 = ~((shr_mem_8_cns_ppown==2'b10));
  assign shr_mem_8_cns_S0_pff = ~((shr_mem_8_acc_rmff==2'b10));
  assign shr_mem_8_mux_6_nl = MUX_s_1_2_2(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_8_and_3_cse_pff);
  assign shr_mem_8_shr_mem_8_or_cse_pff = (shr_mem_8_mux_6_nl) | (~((shr_mem_8_cns_S0_pff
      & (~ shr_mem_8_xor_rmff)) | shr_mem_8_and_3_cse_pff));
  assign shr_mem_8_cns_csb_n_shi0 = shr_mem_8_shr_mem_8_or_cse_pff;
  assign shr_mem_8_cns_dinb_shi0 = MUX_v_64_2_2(dout_8_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_8_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_8_and_3_cse_pff);
  assign shr_mem_8_cns_addra_shi1 = shr_mem_8_shr_mem_8_mux_2_cse_pff;
  assign shr_mem_8_and_5_cse_pff = shr_mem_8_cns_S1_pff & shr_mem_8_xor_1_rmff;
  assign shr_mem_8_shr_mem_8_mux_2_cse_pff = MUX_v_7_2_2(dout_8_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_8_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_8_and_5_cse_pff);
  assign shr_mem_8_cns_addrb_shi1 = shr_mem_8_shr_mem_8_mux_2_cse_pff;
  assign shr_mem_8_cns_csa_n_shi1 = shr_mem_8_shr_mem_8_or_1_cse_pff;
  assign shr_mem_8_mux_7_nl = MUX_s_1_2_2(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_8_and_5_cse_pff);
  assign shr_mem_8_shr_mem_8_or_1_cse_pff = (shr_mem_8_mux_7_nl) | (~((shr_mem_8_cns_S0_pff
      & shr_mem_8_xor_rmff) | shr_mem_8_and_5_cse_pff));
  assign shr_mem_8_cns_csb_n_shi1 = shr_mem_8_shr_mem_8_or_1_cse_pff;
  assign shr_mem_8_cns_dinb_shi1 = MUX_v_64_2_2(dout_8_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_8_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_8_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_8_cns_ppidx <= 1'b0;
      shr_mem_8_cns_ppown <= 2'b0;
      shr_mem_8_cns_ppidx_1 <= 1'b0;
      shr_mem_8_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_8_cns_ppidx <= shr_mem_8_xor_rmff;
      shr_mem_8_cns_ppown <= shr_mem_8_acc_rmff;
      shr_mem_8_cns_ppidx_1 <= shr_mem_8_xor_1_rmff;
      shr_mem_8_cns_ppown_1 <= shr_mem_8_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeaIgYu_7_cns_bctl
// ------------------------------------------------------------------


module double_buffeaIgYu_7_cns_bctl (
  clk, rst, dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_7_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_7_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_7_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_7_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_7_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_7_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_7_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_7_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_7_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_7_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_7_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_7_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_7_cns_S0, shr_mem_7_cns_R0, shr_mem_7_cns_S1, shr_mem_7_cns_R1, shr_mem_7_cns_addra_shi0,
      shr_mem_7_cns_addra_shi1, shr_mem_7_cns_addrb_shi0, shr_mem_7_cns_addrb_shi1,
      shr_mem_7_cns_csa_n_shi0, shr_mem_7_cns_csa_n_shi1, shr_mem_7_cns_csb_n_shi0,
      shr_mem_7_cns_csb_n_shi1, shr_mem_7_cns_dinb_shi0, shr_mem_7_cns_dinb_shi1,
      shr_mem_7_cns_douta_sho0, shr_mem_7_cns_douta_sho1, shr_mem_7_cns_S1_pff, din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_7_cns_S0_pff
);
  input clk;
  input rst;
  input dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_7_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_7_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_7_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_7_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_7_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_7_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_7_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_7_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_7_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_7_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_7_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_7_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_7_cns_S0;
  input shr_mem_7_cns_R0;
  output shr_mem_7_cns_S1;
  input shr_mem_7_cns_R1;
  output [6:0] shr_mem_7_cns_addra_shi0;
  output [6:0] shr_mem_7_cns_addra_shi1;
  output [6:0] shr_mem_7_cns_addrb_shi0;
  output [6:0] shr_mem_7_cns_addrb_shi1;
  output shr_mem_7_cns_csa_n_shi0;
  output shr_mem_7_cns_csa_n_shi1;
  output shr_mem_7_cns_csb_n_shi0;
  output shr_mem_7_cns_csb_n_shi1;
  output [63:0] shr_mem_7_cns_dinb_shi0;
  output [63:0] shr_mem_7_cns_dinb_shi1;
  input [63:0] shr_mem_7_cns_douta_sho0;
  input [63:0] shr_mem_7_cns_douta_sho1;
  output shr_mem_7_cns_S1_pff;
  input din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_7_cns_S0_pff;


  // Interconnect Declarations
  reg dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_7_cns_PC0;
  reg shr_mem_7_cns_ppidx;
  reg [1:0] shr_mem_7_cns_ppown;
  wire shr_mem_7_cns_PC1;
  reg shr_mem_7_cns_ppidx_1;
  reg [1:0] shr_mem_7_cns_ppown_1;
  wire [6:0] shr_mem_7_shr_mem_7_mux_3_cse_pff;
  wire shr_mem_7_and_3_cse_pff;
  wire [1:0] shr_mem_7_acc_1_rmff;
  wire [3:0] nl_shr_mem_7_acc_1_rmff;
  wire shr_mem_7_xor_1_rmff;
  wire shr_mem_7_shr_mem_7_or_cse_pff;
  wire [1:0] shr_mem_7_acc_rmff;
  wire [3:0] nl_shr_mem_7_acc_rmff;
  wire shr_mem_7_xor_rmff;
  wire [6:0] shr_mem_7_shr_mem_7_mux_2_cse_pff;
  wire shr_mem_7_and_5_cse_pff;
  wire shr_mem_7_shr_mem_7_or_1_cse_pff;

  wire[0:0] shr_mem_7_mux_6_nl;
  wire[0:0] shr_mem_7_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_7_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_7_cns_R0;
  assign din_7_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_7_cns_R1;
  assign shr_mem_7_xor_rmff = shr_mem_7_cns_ppidx ^ shr_mem_7_cns_PC0;
  assign nl_shr_mem_7_acc_rmff = shr_mem_7_cns_ppown + conv_u2u_1_2(shr_mem_7_cns_PC0)
      + conv_s2u_1_2(shr_mem_7_cns_PC1);
  assign shr_mem_7_acc_rmff = nl_shr_mem_7_acc_rmff[1:0];
  assign shr_mem_7_cns_PC0 = shr_mem_7_cns_S0 & dout_7_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_7_xor_1_rmff = shr_mem_7_cns_ppidx_1 ^ shr_mem_7_cns_PC1;
  assign nl_shr_mem_7_acc_1_rmff = shr_mem_7_cns_ppown_1 + conv_u2u_1_2(shr_mem_7_cns_PC1)
      + conv_s2u_1_2(shr_mem_7_cns_PC0);
  assign shr_mem_7_acc_1_rmff = nl_shr_mem_7_acc_1_rmff[1:0];
  assign shr_mem_7_cns_PC1 = shr_mem_7_cns_S1 & din_7_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_7_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_7_cns_douta_sho0,
      shr_mem_7_cns_douta_sho1, shr_mem_7_cns_ppidx);
  assign din_7_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_7_cns_douta_sho0,
      shr_mem_7_cns_douta_sho1, shr_mem_7_cns_ppidx_1);
  assign shr_mem_7_cns_addra_shi0 = shr_mem_7_shr_mem_7_mux_3_cse_pff;
  assign shr_mem_7_cns_S1 = (shr_mem_7_cns_ppown_1!=2'b00);
  assign shr_mem_7_cns_S1_pff = (shr_mem_7_acc_1_rmff!=2'b00);
  assign shr_mem_7_and_3_cse_pff = shr_mem_7_cns_S1_pff & (~ shr_mem_7_xor_1_rmff);
  assign shr_mem_7_shr_mem_7_mux_3_cse_pff = MUX_v_7_2_2(dout_7_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_7_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_7_and_3_cse_pff);
  assign shr_mem_7_cns_addrb_shi0 = shr_mem_7_shr_mem_7_mux_3_cse_pff;
  assign shr_mem_7_cns_csa_n_shi0 = shr_mem_7_shr_mem_7_or_cse_pff;
  assign din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff = din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff = dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_7_cns_S0 = ~((shr_mem_7_cns_ppown==2'b10));
  assign shr_mem_7_cns_S0_pff = ~((shr_mem_7_acc_rmff==2'b10));
  assign shr_mem_7_mux_6_nl = MUX_s_1_2_2(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_7_and_3_cse_pff);
  assign shr_mem_7_shr_mem_7_or_cse_pff = (shr_mem_7_mux_6_nl) | (~((shr_mem_7_cns_S0_pff
      & (~ shr_mem_7_xor_rmff)) | shr_mem_7_and_3_cse_pff));
  assign shr_mem_7_cns_csb_n_shi0 = shr_mem_7_shr_mem_7_or_cse_pff;
  assign shr_mem_7_cns_dinb_shi0 = MUX_v_64_2_2(dout_7_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_7_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_7_and_3_cse_pff);
  assign shr_mem_7_cns_addra_shi1 = shr_mem_7_shr_mem_7_mux_2_cse_pff;
  assign shr_mem_7_and_5_cse_pff = shr_mem_7_cns_S1_pff & shr_mem_7_xor_1_rmff;
  assign shr_mem_7_shr_mem_7_mux_2_cse_pff = MUX_v_7_2_2(dout_7_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_7_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_7_and_5_cse_pff);
  assign shr_mem_7_cns_addrb_shi1 = shr_mem_7_shr_mem_7_mux_2_cse_pff;
  assign shr_mem_7_cns_csa_n_shi1 = shr_mem_7_shr_mem_7_or_1_cse_pff;
  assign shr_mem_7_mux_7_nl = MUX_s_1_2_2(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_7_and_5_cse_pff);
  assign shr_mem_7_shr_mem_7_or_1_cse_pff = (shr_mem_7_mux_7_nl) | (~((shr_mem_7_cns_S0_pff
      & shr_mem_7_xor_rmff) | shr_mem_7_and_5_cse_pff));
  assign shr_mem_7_cns_csb_n_shi1 = shr_mem_7_shr_mem_7_or_1_cse_pff;
  assign shr_mem_7_cns_dinb_shi1 = MUX_v_64_2_2(dout_7_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_7_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_7_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_7_cns_ppidx <= 1'b0;
      shr_mem_7_cns_ppown <= 2'b0;
      shr_mem_7_cns_ppidx_1 <= 1'b0;
      shr_mem_7_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_7_cns_ppidx <= shr_mem_7_xor_rmff;
      shr_mem_7_cns_ppown <= shr_mem_7_acc_rmff;
      shr_mem_7_cns_ppidx_1 <= shr_mem_7_xor_1_rmff;
      shr_mem_7_cns_ppown_1 <= shr_mem_7_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeaIgYu_6_cns_bctl
// ------------------------------------------------------------------


module double_buffeaIgYu_6_cns_bctl (
  clk, rst, dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_6_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_6_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_6_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_6_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_6_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_6_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_6_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_6_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_6_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_6_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_6_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_6_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_6_cns_S0, shr_mem_6_cns_R0, shr_mem_6_cns_S1, shr_mem_6_cns_R1, shr_mem_6_cns_addra_shi0,
      shr_mem_6_cns_addra_shi1, shr_mem_6_cns_addrb_shi0, shr_mem_6_cns_addrb_shi1,
      shr_mem_6_cns_csa_n_shi0, shr_mem_6_cns_csa_n_shi1, shr_mem_6_cns_csb_n_shi0,
      shr_mem_6_cns_csb_n_shi1, shr_mem_6_cns_dinb_shi0, shr_mem_6_cns_dinb_shi1,
      shr_mem_6_cns_douta_sho0, shr_mem_6_cns_douta_sho1, shr_mem_6_cns_S1_pff, din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_6_cns_S0_pff
);
  input clk;
  input rst;
  input dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_6_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_6_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_6_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_6_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_6_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_6_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_6_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_6_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_6_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_6_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_6_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_6_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_6_cns_S0;
  input shr_mem_6_cns_R0;
  output shr_mem_6_cns_S1;
  input shr_mem_6_cns_R1;
  output [6:0] shr_mem_6_cns_addra_shi0;
  output [6:0] shr_mem_6_cns_addra_shi1;
  output [6:0] shr_mem_6_cns_addrb_shi0;
  output [6:0] shr_mem_6_cns_addrb_shi1;
  output shr_mem_6_cns_csa_n_shi0;
  output shr_mem_6_cns_csa_n_shi1;
  output shr_mem_6_cns_csb_n_shi0;
  output shr_mem_6_cns_csb_n_shi1;
  output [63:0] shr_mem_6_cns_dinb_shi0;
  output [63:0] shr_mem_6_cns_dinb_shi1;
  input [63:0] shr_mem_6_cns_douta_sho0;
  input [63:0] shr_mem_6_cns_douta_sho1;
  output shr_mem_6_cns_S1_pff;
  input din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_6_cns_S0_pff;


  // Interconnect Declarations
  reg dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_6_cns_PC0;
  reg shr_mem_6_cns_ppidx;
  reg [1:0] shr_mem_6_cns_ppown;
  wire shr_mem_6_cns_PC1;
  reg shr_mem_6_cns_ppidx_1;
  reg [1:0] shr_mem_6_cns_ppown_1;
  wire [6:0] shr_mem_6_shr_mem_6_mux_3_cse_pff;
  wire shr_mem_6_and_3_cse_pff;
  wire [1:0] shr_mem_6_acc_1_rmff;
  wire [3:0] nl_shr_mem_6_acc_1_rmff;
  wire shr_mem_6_xor_1_rmff;
  wire shr_mem_6_shr_mem_6_or_cse_pff;
  wire [1:0] shr_mem_6_acc_rmff;
  wire [3:0] nl_shr_mem_6_acc_rmff;
  wire shr_mem_6_xor_rmff;
  wire [6:0] shr_mem_6_shr_mem_6_mux_2_cse_pff;
  wire shr_mem_6_and_5_cse_pff;
  wire shr_mem_6_shr_mem_6_or_1_cse_pff;

  wire[0:0] shr_mem_6_mux_6_nl;
  wire[0:0] shr_mem_6_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_6_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_6_cns_R0;
  assign din_6_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_6_cns_R1;
  assign shr_mem_6_xor_rmff = shr_mem_6_cns_ppidx ^ shr_mem_6_cns_PC0;
  assign nl_shr_mem_6_acc_rmff = shr_mem_6_cns_ppown + conv_u2u_1_2(shr_mem_6_cns_PC0)
      + conv_s2u_1_2(shr_mem_6_cns_PC1);
  assign shr_mem_6_acc_rmff = nl_shr_mem_6_acc_rmff[1:0];
  assign shr_mem_6_cns_PC0 = shr_mem_6_cns_S0 & dout_6_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_6_xor_1_rmff = shr_mem_6_cns_ppidx_1 ^ shr_mem_6_cns_PC1;
  assign nl_shr_mem_6_acc_1_rmff = shr_mem_6_cns_ppown_1 + conv_u2u_1_2(shr_mem_6_cns_PC1)
      + conv_s2u_1_2(shr_mem_6_cns_PC0);
  assign shr_mem_6_acc_1_rmff = nl_shr_mem_6_acc_1_rmff[1:0];
  assign shr_mem_6_cns_PC1 = shr_mem_6_cns_S1 & din_6_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_6_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_6_cns_douta_sho0,
      shr_mem_6_cns_douta_sho1, shr_mem_6_cns_ppidx);
  assign din_6_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_6_cns_douta_sho0,
      shr_mem_6_cns_douta_sho1, shr_mem_6_cns_ppidx_1);
  assign shr_mem_6_cns_addra_shi0 = shr_mem_6_shr_mem_6_mux_3_cse_pff;
  assign shr_mem_6_cns_S1 = (shr_mem_6_cns_ppown_1!=2'b00);
  assign shr_mem_6_cns_S1_pff = (shr_mem_6_acc_1_rmff!=2'b00);
  assign shr_mem_6_and_3_cse_pff = shr_mem_6_cns_S1_pff & (~ shr_mem_6_xor_1_rmff);
  assign shr_mem_6_shr_mem_6_mux_3_cse_pff = MUX_v_7_2_2(dout_6_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_6_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_6_and_3_cse_pff);
  assign shr_mem_6_cns_addrb_shi0 = shr_mem_6_shr_mem_6_mux_3_cse_pff;
  assign shr_mem_6_cns_csa_n_shi0 = shr_mem_6_shr_mem_6_or_cse_pff;
  assign din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff = din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff = dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_6_cns_S0 = ~((shr_mem_6_cns_ppown==2'b10));
  assign shr_mem_6_cns_S0_pff = ~((shr_mem_6_acc_rmff==2'b10));
  assign shr_mem_6_mux_6_nl = MUX_s_1_2_2(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_6_and_3_cse_pff);
  assign shr_mem_6_shr_mem_6_or_cse_pff = (shr_mem_6_mux_6_nl) | (~((shr_mem_6_cns_S0_pff
      & (~ shr_mem_6_xor_rmff)) | shr_mem_6_and_3_cse_pff));
  assign shr_mem_6_cns_csb_n_shi0 = shr_mem_6_shr_mem_6_or_cse_pff;
  assign shr_mem_6_cns_dinb_shi0 = MUX_v_64_2_2(dout_6_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_6_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_6_and_3_cse_pff);
  assign shr_mem_6_cns_addra_shi1 = shr_mem_6_shr_mem_6_mux_2_cse_pff;
  assign shr_mem_6_and_5_cse_pff = shr_mem_6_cns_S1_pff & shr_mem_6_xor_1_rmff;
  assign shr_mem_6_shr_mem_6_mux_2_cse_pff = MUX_v_7_2_2(dout_6_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_6_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_6_and_5_cse_pff);
  assign shr_mem_6_cns_addrb_shi1 = shr_mem_6_shr_mem_6_mux_2_cse_pff;
  assign shr_mem_6_cns_csa_n_shi1 = shr_mem_6_shr_mem_6_or_1_cse_pff;
  assign shr_mem_6_mux_7_nl = MUX_s_1_2_2(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_6_and_5_cse_pff);
  assign shr_mem_6_shr_mem_6_or_1_cse_pff = (shr_mem_6_mux_7_nl) | (~((shr_mem_6_cns_S0_pff
      & shr_mem_6_xor_rmff) | shr_mem_6_and_5_cse_pff));
  assign shr_mem_6_cns_csb_n_shi1 = shr_mem_6_shr_mem_6_or_1_cse_pff;
  assign shr_mem_6_cns_dinb_shi1 = MUX_v_64_2_2(dout_6_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_6_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_6_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_6_cns_ppidx <= 1'b0;
      shr_mem_6_cns_ppown <= 2'b0;
      shr_mem_6_cns_ppidx_1 <= 1'b0;
      shr_mem_6_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_6_cns_ppidx <= shr_mem_6_xor_rmff;
      shr_mem_6_cns_ppown <= shr_mem_6_acc_rmff;
      shr_mem_6_cns_ppidx_1 <= shr_mem_6_xor_1_rmff;
      shr_mem_6_cns_ppown_1 <= shr_mem_6_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeaIgYu_5_cns_bctl
// ------------------------------------------------------------------


module double_buffeaIgYu_5_cns_bctl (
  clk, rst, dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_5_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_5_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_5_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_5_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_5_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_5_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_5_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_5_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_5_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_5_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_5_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_5_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_5_cns_S0, shr_mem_5_cns_R0, shr_mem_5_cns_S1, shr_mem_5_cns_R1, shr_mem_5_cns_addra_shi0,
      shr_mem_5_cns_addra_shi1, shr_mem_5_cns_addrb_shi0, shr_mem_5_cns_addrb_shi1,
      shr_mem_5_cns_csa_n_shi0, shr_mem_5_cns_csa_n_shi1, shr_mem_5_cns_csb_n_shi0,
      shr_mem_5_cns_csb_n_shi1, shr_mem_5_cns_dinb_shi0, shr_mem_5_cns_dinb_shi1,
      shr_mem_5_cns_douta_sho0, shr_mem_5_cns_douta_sho1, shr_mem_5_cns_S1_pff, din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_5_cns_S0_pff
);
  input clk;
  input rst;
  input dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_5_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_5_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_5_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_5_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_5_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_5_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_5_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_5_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_5_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_5_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_5_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_5_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_5_cns_S0;
  input shr_mem_5_cns_R0;
  output shr_mem_5_cns_S1;
  input shr_mem_5_cns_R1;
  output [6:0] shr_mem_5_cns_addra_shi0;
  output [6:0] shr_mem_5_cns_addra_shi1;
  output [6:0] shr_mem_5_cns_addrb_shi0;
  output [6:0] shr_mem_5_cns_addrb_shi1;
  output shr_mem_5_cns_csa_n_shi0;
  output shr_mem_5_cns_csa_n_shi1;
  output shr_mem_5_cns_csb_n_shi0;
  output shr_mem_5_cns_csb_n_shi1;
  output [63:0] shr_mem_5_cns_dinb_shi0;
  output [63:0] shr_mem_5_cns_dinb_shi1;
  input [63:0] shr_mem_5_cns_douta_sho0;
  input [63:0] shr_mem_5_cns_douta_sho1;
  output shr_mem_5_cns_S1_pff;
  input din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_5_cns_S0_pff;


  // Interconnect Declarations
  reg dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_5_cns_PC0;
  reg shr_mem_5_cns_ppidx;
  reg [1:0] shr_mem_5_cns_ppown;
  wire shr_mem_5_cns_PC1;
  reg shr_mem_5_cns_ppidx_1;
  reg [1:0] shr_mem_5_cns_ppown_1;
  wire [6:0] shr_mem_5_shr_mem_5_mux_3_cse_pff;
  wire shr_mem_5_and_3_cse_pff;
  wire [1:0] shr_mem_5_acc_1_rmff;
  wire [3:0] nl_shr_mem_5_acc_1_rmff;
  wire shr_mem_5_xor_1_rmff;
  wire shr_mem_5_shr_mem_5_or_cse_pff;
  wire [1:0] shr_mem_5_acc_rmff;
  wire [3:0] nl_shr_mem_5_acc_rmff;
  wire shr_mem_5_xor_rmff;
  wire [6:0] shr_mem_5_shr_mem_5_mux_2_cse_pff;
  wire shr_mem_5_and_5_cse_pff;
  wire shr_mem_5_shr_mem_5_or_1_cse_pff;

  wire[0:0] shr_mem_5_mux_6_nl;
  wire[0:0] shr_mem_5_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_5_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_5_cns_R0;
  assign din_5_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_5_cns_R1;
  assign shr_mem_5_xor_rmff = shr_mem_5_cns_ppidx ^ shr_mem_5_cns_PC0;
  assign nl_shr_mem_5_acc_rmff = shr_mem_5_cns_ppown + conv_u2u_1_2(shr_mem_5_cns_PC0)
      + conv_s2u_1_2(shr_mem_5_cns_PC1);
  assign shr_mem_5_acc_rmff = nl_shr_mem_5_acc_rmff[1:0];
  assign shr_mem_5_cns_PC0 = shr_mem_5_cns_S0 & dout_5_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_5_xor_1_rmff = shr_mem_5_cns_ppidx_1 ^ shr_mem_5_cns_PC1;
  assign nl_shr_mem_5_acc_1_rmff = shr_mem_5_cns_ppown_1 + conv_u2u_1_2(shr_mem_5_cns_PC1)
      + conv_s2u_1_2(shr_mem_5_cns_PC0);
  assign shr_mem_5_acc_1_rmff = nl_shr_mem_5_acc_1_rmff[1:0];
  assign shr_mem_5_cns_PC1 = shr_mem_5_cns_S1 & din_5_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_5_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_5_cns_douta_sho0,
      shr_mem_5_cns_douta_sho1, shr_mem_5_cns_ppidx);
  assign din_5_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_5_cns_douta_sho0,
      shr_mem_5_cns_douta_sho1, shr_mem_5_cns_ppidx_1);
  assign shr_mem_5_cns_addra_shi0 = shr_mem_5_shr_mem_5_mux_3_cse_pff;
  assign shr_mem_5_cns_S1 = (shr_mem_5_cns_ppown_1!=2'b00);
  assign shr_mem_5_cns_S1_pff = (shr_mem_5_acc_1_rmff!=2'b00);
  assign shr_mem_5_and_3_cse_pff = shr_mem_5_cns_S1_pff & (~ shr_mem_5_xor_1_rmff);
  assign shr_mem_5_shr_mem_5_mux_3_cse_pff = MUX_v_7_2_2(dout_5_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_5_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_5_and_3_cse_pff);
  assign shr_mem_5_cns_addrb_shi0 = shr_mem_5_shr_mem_5_mux_3_cse_pff;
  assign shr_mem_5_cns_csa_n_shi0 = shr_mem_5_shr_mem_5_or_cse_pff;
  assign din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff = din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff = dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_5_cns_S0 = ~((shr_mem_5_cns_ppown==2'b10));
  assign shr_mem_5_cns_S0_pff = ~((shr_mem_5_acc_rmff==2'b10));
  assign shr_mem_5_mux_6_nl = MUX_s_1_2_2(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_5_and_3_cse_pff);
  assign shr_mem_5_shr_mem_5_or_cse_pff = (shr_mem_5_mux_6_nl) | (~((shr_mem_5_cns_S0_pff
      & (~ shr_mem_5_xor_rmff)) | shr_mem_5_and_3_cse_pff));
  assign shr_mem_5_cns_csb_n_shi0 = shr_mem_5_shr_mem_5_or_cse_pff;
  assign shr_mem_5_cns_dinb_shi0 = MUX_v_64_2_2(dout_5_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_5_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_5_and_3_cse_pff);
  assign shr_mem_5_cns_addra_shi1 = shr_mem_5_shr_mem_5_mux_2_cse_pff;
  assign shr_mem_5_and_5_cse_pff = shr_mem_5_cns_S1_pff & shr_mem_5_xor_1_rmff;
  assign shr_mem_5_shr_mem_5_mux_2_cse_pff = MUX_v_7_2_2(dout_5_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_5_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_5_and_5_cse_pff);
  assign shr_mem_5_cns_addrb_shi1 = shr_mem_5_shr_mem_5_mux_2_cse_pff;
  assign shr_mem_5_cns_csa_n_shi1 = shr_mem_5_shr_mem_5_or_1_cse_pff;
  assign shr_mem_5_mux_7_nl = MUX_s_1_2_2(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_5_and_5_cse_pff);
  assign shr_mem_5_shr_mem_5_or_1_cse_pff = (shr_mem_5_mux_7_nl) | (~((shr_mem_5_cns_S0_pff
      & shr_mem_5_xor_rmff) | shr_mem_5_and_5_cse_pff));
  assign shr_mem_5_cns_csb_n_shi1 = shr_mem_5_shr_mem_5_or_1_cse_pff;
  assign shr_mem_5_cns_dinb_shi1 = MUX_v_64_2_2(dout_5_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_5_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_5_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_5_cns_ppidx <= 1'b0;
      shr_mem_5_cns_ppown <= 2'b0;
      shr_mem_5_cns_ppidx_1 <= 1'b0;
      shr_mem_5_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_5_cns_ppidx <= shr_mem_5_xor_rmff;
      shr_mem_5_cns_ppown <= shr_mem_5_acc_rmff;
      shr_mem_5_cns_ppidx_1 <= shr_mem_5_xor_1_rmff;
      shr_mem_5_cns_ppown_1 <= shr_mem_5_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeaIgYu_4_cns_bctl
// ------------------------------------------------------------------


module double_buffeaIgYu_4_cns_bctl (
  clk, rst, dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_4_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_4_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_4_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_4_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_4_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_4_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_4_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_4_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_4_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_4_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_4_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_4_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_4_cns_S0, shr_mem_4_cns_R0, shr_mem_4_cns_S1, shr_mem_4_cns_R1, shr_mem_4_cns_addra_shi0,
      shr_mem_4_cns_addra_shi1, shr_mem_4_cns_addrb_shi0, shr_mem_4_cns_addrb_shi1,
      shr_mem_4_cns_csa_n_shi0, shr_mem_4_cns_csa_n_shi1, shr_mem_4_cns_csb_n_shi0,
      shr_mem_4_cns_csb_n_shi1, shr_mem_4_cns_dinb_shi0, shr_mem_4_cns_dinb_shi1,
      shr_mem_4_cns_douta_sho0, shr_mem_4_cns_douta_sho1, shr_mem_4_cns_S1_pff, din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_4_cns_S0_pff
);
  input clk;
  input rst;
  input dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_4_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_4_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_4_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_4_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_4_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_4_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_4_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_4_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_4_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_4_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_4_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_4_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_4_cns_S0;
  input shr_mem_4_cns_R0;
  output shr_mem_4_cns_S1;
  input shr_mem_4_cns_R1;
  output [6:0] shr_mem_4_cns_addra_shi0;
  output [6:0] shr_mem_4_cns_addra_shi1;
  output [6:0] shr_mem_4_cns_addrb_shi0;
  output [6:0] shr_mem_4_cns_addrb_shi1;
  output shr_mem_4_cns_csa_n_shi0;
  output shr_mem_4_cns_csa_n_shi1;
  output shr_mem_4_cns_csb_n_shi0;
  output shr_mem_4_cns_csb_n_shi1;
  output [63:0] shr_mem_4_cns_dinb_shi0;
  output [63:0] shr_mem_4_cns_dinb_shi1;
  input [63:0] shr_mem_4_cns_douta_sho0;
  input [63:0] shr_mem_4_cns_douta_sho1;
  output shr_mem_4_cns_S1_pff;
  input din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_4_cns_S0_pff;


  // Interconnect Declarations
  reg dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_4_cns_PC0;
  reg shr_mem_4_cns_ppidx;
  reg [1:0] shr_mem_4_cns_ppown;
  wire shr_mem_4_cns_PC1;
  reg shr_mem_4_cns_ppidx_1;
  reg [1:0] shr_mem_4_cns_ppown_1;
  wire [6:0] shr_mem_4_shr_mem_4_mux_3_cse_pff;
  wire shr_mem_4_and_3_cse_pff;
  wire [1:0] shr_mem_4_acc_1_rmff;
  wire [3:0] nl_shr_mem_4_acc_1_rmff;
  wire shr_mem_4_xor_1_rmff;
  wire shr_mem_4_shr_mem_4_or_cse_pff;
  wire [1:0] shr_mem_4_acc_rmff;
  wire [3:0] nl_shr_mem_4_acc_rmff;
  wire shr_mem_4_xor_rmff;
  wire [6:0] shr_mem_4_shr_mem_4_mux_2_cse_pff;
  wire shr_mem_4_and_5_cse_pff;
  wire shr_mem_4_shr_mem_4_or_1_cse_pff;

  wire[0:0] shr_mem_4_mux_6_nl;
  wire[0:0] shr_mem_4_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_4_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_4_cns_R0;
  assign din_4_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_4_cns_R1;
  assign shr_mem_4_xor_rmff = shr_mem_4_cns_ppidx ^ shr_mem_4_cns_PC0;
  assign nl_shr_mem_4_acc_rmff = shr_mem_4_cns_ppown + conv_u2u_1_2(shr_mem_4_cns_PC0)
      + conv_s2u_1_2(shr_mem_4_cns_PC1);
  assign shr_mem_4_acc_rmff = nl_shr_mem_4_acc_rmff[1:0];
  assign shr_mem_4_cns_PC0 = shr_mem_4_cns_S0 & dout_4_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_4_xor_1_rmff = shr_mem_4_cns_ppidx_1 ^ shr_mem_4_cns_PC1;
  assign nl_shr_mem_4_acc_1_rmff = shr_mem_4_cns_ppown_1 + conv_u2u_1_2(shr_mem_4_cns_PC1)
      + conv_s2u_1_2(shr_mem_4_cns_PC0);
  assign shr_mem_4_acc_1_rmff = nl_shr_mem_4_acc_1_rmff[1:0];
  assign shr_mem_4_cns_PC1 = shr_mem_4_cns_S1 & din_4_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_4_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_4_cns_douta_sho0,
      shr_mem_4_cns_douta_sho1, shr_mem_4_cns_ppidx);
  assign din_4_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_4_cns_douta_sho0,
      shr_mem_4_cns_douta_sho1, shr_mem_4_cns_ppidx_1);
  assign shr_mem_4_cns_addra_shi0 = shr_mem_4_shr_mem_4_mux_3_cse_pff;
  assign shr_mem_4_cns_S1 = (shr_mem_4_cns_ppown_1!=2'b00);
  assign shr_mem_4_cns_S1_pff = (shr_mem_4_acc_1_rmff!=2'b00);
  assign shr_mem_4_and_3_cse_pff = shr_mem_4_cns_S1_pff & (~ shr_mem_4_xor_1_rmff);
  assign shr_mem_4_shr_mem_4_mux_3_cse_pff = MUX_v_7_2_2(dout_4_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_4_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_4_and_3_cse_pff);
  assign shr_mem_4_cns_addrb_shi0 = shr_mem_4_shr_mem_4_mux_3_cse_pff;
  assign shr_mem_4_cns_csa_n_shi0 = shr_mem_4_shr_mem_4_or_cse_pff;
  assign din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff = din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff = dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_4_cns_S0 = ~((shr_mem_4_cns_ppown==2'b10));
  assign shr_mem_4_cns_S0_pff = ~((shr_mem_4_acc_rmff==2'b10));
  assign shr_mem_4_mux_6_nl = MUX_s_1_2_2(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_4_and_3_cse_pff);
  assign shr_mem_4_shr_mem_4_or_cse_pff = (shr_mem_4_mux_6_nl) | (~((shr_mem_4_cns_S0_pff
      & (~ shr_mem_4_xor_rmff)) | shr_mem_4_and_3_cse_pff));
  assign shr_mem_4_cns_csb_n_shi0 = shr_mem_4_shr_mem_4_or_cse_pff;
  assign shr_mem_4_cns_dinb_shi0 = MUX_v_64_2_2(dout_4_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_4_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_4_and_3_cse_pff);
  assign shr_mem_4_cns_addra_shi1 = shr_mem_4_shr_mem_4_mux_2_cse_pff;
  assign shr_mem_4_and_5_cse_pff = shr_mem_4_cns_S1_pff & shr_mem_4_xor_1_rmff;
  assign shr_mem_4_shr_mem_4_mux_2_cse_pff = MUX_v_7_2_2(dout_4_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_4_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_4_and_5_cse_pff);
  assign shr_mem_4_cns_addrb_shi1 = shr_mem_4_shr_mem_4_mux_2_cse_pff;
  assign shr_mem_4_cns_csa_n_shi1 = shr_mem_4_shr_mem_4_or_1_cse_pff;
  assign shr_mem_4_mux_7_nl = MUX_s_1_2_2(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_4_and_5_cse_pff);
  assign shr_mem_4_shr_mem_4_or_1_cse_pff = (shr_mem_4_mux_7_nl) | (~((shr_mem_4_cns_S0_pff
      & shr_mem_4_xor_rmff) | shr_mem_4_and_5_cse_pff));
  assign shr_mem_4_cns_csb_n_shi1 = shr_mem_4_shr_mem_4_or_1_cse_pff;
  assign shr_mem_4_cns_dinb_shi1 = MUX_v_64_2_2(dout_4_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_4_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_4_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_4_cns_ppidx <= 1'b0;
      shr_mem_4_cns_ppown <= 2'b0;
      shr_mem_4_cns_ppidx_1 <= 1'b0;
      shr_mem_4_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_4_cns_ppidx <= shr_mem_4_xor_rmff;
      shr_mem_4_cns_ppown <= shr_mem_4_acc_rmff;
      shr_mem_4_cns_ppidx_1 <= shr_mem_4_xor_1_rmff;
      shr_mem_4_cns_ppown_1 <= shr_mem_4_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeaIgYu_3_cns_bctl
// ------------------------------------------------------------------


module double_buffeaIgYu_3_cns_bctl (
  clk, rst, dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_3_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_3_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_3_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_3_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_3_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_3_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_3_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_3_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_3_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_3_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_3_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_3_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_3_cns_S0, shr_mem_3_cns_R0, shr_mem_3_cns_S1, shr_mem_3_cns_R1, shr_mem_3_cns_addra_shi0,
      shr_mem_3_cns_addra_shi1, shr_mem_3_cns_addrb_shi0, shr_mem_3_cns_addrb_shi1,
      shr_mem_3_cns_csa_n_shi0, shr_mem_3_cns_csa_n_shi1, shr_mem_3_cns_csb_n_shi0,
      shr_mem_3_cns_csb_n_shi1, shr_mem_3_cns_dinb_shi0, shr_mem_3_cns_dinb_shi1,
      shr_mem_3_cns_douta_sho0, shr_mem_3_cns_douta_sho1, shr_mem_3_cns_S1_pff, din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_3_cns_S0_pff
);
  input clk;
  input rst;
  input dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_3_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_3_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_3_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_3_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_3_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_3_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_3_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_3_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_3_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_3_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_3_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_3_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_3_cns_S0;
  input shr_mem_3_cns_R0;
  output shr_mem_3_cns_S1;
  input shr_mem_3_cns_R1;
  output [6:0] shr_mem_3_cns_addra_shi0;
  output [6:0] shr_mem_3_cns_addra_shi1;
  output [6:0] shr_mem_3_cns_addrb_shi0;
  output [6:0] shr_mem_3_cns_addrb_shi1;
  output shr_mem_3_cns_csa_n_shi0;
  output shr_mem_3_cns_csa_n_shi1;
  output shr_mem_3_cns_csb_n_shi0;
  output shr_mem_3_cns_csb_n_shi1;
  output [63:0] shr_mem_3_cns_dinb_shi0;
  output [63:0] shr_mem_3_cns_dinb_shi1;
  input [63:0] shr_mem_3_cns_douta_sho0;
  input [63:0] shr_mem_3_cns_douta_sho1;
  output shr_mem_3_cns_S1_pff;
  input din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_3_cns_S0_pff;


  // Interconnect Declarations
  reg dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_3_cns_PC0;
  reg shr_mem_3_cns_ppidx;
  reg [1:0] shr_mem_3_cns_ppown;
  wire shr_mem_3_cns_PC1;
  reg shr_mem_3_cns_ppidx_1;
  reg [1:0] shr_mem_3_cns_ppown_1;
  wire [6:0] shr_mem_3_shr_mem_3_mux_3_cse_pff;
  wire shr_mem_3_and_3_cse_pff;
  wire [1:0] shr_mem_3_acc_1_rmff;
  wire [3:0] nl_shr_mem_3_acc_1_rmff;
  wire shr_mem_3_xor_1_rmff;
  wire shr_mem_3_shr_mem_3_or_cse_pff;
  wire [1:0] shr_mem_3_acc_rmff;
  wire [3:0] nl_shr_mem_3_acc_rmff;
  wire shr_mem_3_xor_rmff;
  wire [6:0] shr_mem_3_shr_mem_3_mux_2_cse_pff;
  wire shr_mem_3_and_5_cse_pff;
  wire shr_mem_3_shr_mem_3_or_1_cse_pff;

  wire[0:0] shr_mem_3_mux_6_nl;
  wire[0:0] shr_mem_3_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_3_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_3_cns_R0;
  assign din_3_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_3_cns_R1;
  assign shr_mem_3_xor_rmff = shr_mem_3_cns_ppidx ^ shr_mem_3_cns_PC0;
  assign nl_shr_mem_3_acc_rmff = shr_mem_3_cns_ppown + conv_u2u_1_2(shr_mem_3_cns_PC0)
      + conv_s2u_1_2(shr_mem_3_cns_PC1);
  assign shr_mem_3_acc_rmff = nl_shr_mem_3_acc_rmff[1:0];
  assign shr_mem_3_cns_PC0 = shr_mem_3_cns_S0 & dout_3_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_3_xor_1_rmff = shr_mem_3_cns_ppidx_1 ^ shr_mem_3_cns_PC1;
  assign nl_shr_mem_3_acc_1_rmff = shr_mem_3_cns_ppown_1 + conv_u2u_1_2(shr_mem_3_cns_PC1)
      + conv_s2u_1_2(shr_mem_3_cns_PC0);
  assign shr_mem_3_acc_1_rmff = nl_shr_mem_3_acc_1_rmff[1:0];
  assign shr_mem_3_cns_PC1 = shr_mem_3_cns_S1 & din_3_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_3_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_3_cns_douta_sho0,
      shr_mem_3_cns_douta_sho1, shr_mem_3_cns_ppidx);
  assign din_3_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_3_cns_douta_sho0,
      shr_mem_3_cns_douta_sho1, shr_mem_3_cns_ppidx_1);
  assign shr_mem_3_cns_addra_shi0 = shr_mem_3_shr_mem_3_mux_3_cse_pff;
  assign shr_mem_3_cns_S1 = (shr_mem_3_cns_ppown_1!=2'b00);
  assign shr_mem_3_cns_S1_pff = (shr_mem_3_acc_1_rmff!=2'b00);
  assign shr_mem_3_and_3_cse_pff = shr_mem_3_cns_S1_pff & (~ shr_mem_3_xor_1_rmff);
  assign shr_mem_3_shr_mem_3_mux_3_cse_pff = MUX_v_7_2_2(dout_3_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_3_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_3_and_3_cse_pff);
  assign shr_mem_3_cns_addrb_shi0 = shr_mem_3_shr_mem_3_mux_3_cse_pff;
  assign shr_mem_3_cns_csa_n_shi0 = shr_mem_3_shr_mem_3_or_cse_pff;
  assign din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff = din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff = dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_3_cns_S0 = ~((shr_mem_3_cns_ppown==2'b10));
  assign shr_mem_3_cns_S0_pff = ~((shr_mem_3_acc_rmff==2'b10));
  assign shr_mem_3_mux_6_nl = MUX_s_1_2_2(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_3_and_3_cse_pff);
  assign shr_mem_3_shr_mem_3_or_cse_pff = (shr_mem_3_mux_6_nl) | (~((shr_mem_3_cns_S0_pff
      & (~ shr_mem_3_xor_rmff)) | shr_mem_3_and_3_cse_pff));
  assign shr_mem_3_cns_csb_n_shi0 = shr_mem_3_shr_mem_3_or_cse_pff;
  assign shr_mem_3_cns_dinb_shi0 = MUX_v_64_2_2(dout_3_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_3_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_3_and_3_cse_pff);
  assign shr_mem_3_cns_addra_shi1 = shr_mem_3_shr_mem_3_mux_2_cse_pff;
  assign shr_mem_3_and_5_cse_pff = shr_mem_3_cns_S1_pff & shr_mem_3_xor_1_rmff;
  assign shr_mem_3_shr_mem_3_mux_2_cse_pff = MUX_v_7_2_2(dout_3_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_3_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_3_and_5_cse_pff);
  assign shr_mem_3_cns_addrb_shi1 = shr_mem_3_shr_mem_3_mux_2_cse_pff;
  assign shr_mem_3_cns_csa_n_shi1 = shr_mem_3_shr_mem_3_or_1_cse_pff;
  assign shr_mem_3_mux_7_nl = MUX_s_1_2_2(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_3_and_5_cse_pff);
  assign shr_mem_3_shr_mem_3_or_1_cse_pff = (shr_mem_3_mux_7_nl) | (~((shr_mem_3_cns_S0_pff
      & shr_mem_3_xor_rmff) | shr_mem_3_and_5_cse_pff));
  assign shr_mem_3_cns_csb_n_shi1 = shr_mem_3_shr_mem_3_or_1_cse_pff;
  assign shr_mem_3_cns_dinb_shi1 = MUX_v_64_2_2(dout_3_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_3_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_3_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_3_cns_ppidx <= 1'b0;
      shr_mem_3_cns_ppown <= 2'b0;
      shr_mem_3_cns_ppidx_1 <= 1'b0;
      shr_mem_3_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_3_cns_ppidx <= shr_mem_3_xor_rmff;
      shr_mem_3_cns_ppown <= shr_mem_3_acc_rmff;
      shr_mem_3_cns_ppidx_1 <= shr_mem_3_xor_1_rmff;
      shr_mem_3_cns_ppown_1 <= shr_mem_3_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeaIgYu_2_cns_bctl
// ------------------------------------------------------------------


module double_buffeaIgYu_2_cns_bctl (
  clk, rst, dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_2_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_2_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_2_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_2_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_2_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_2_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_2_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_2_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_2_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_2_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_2_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_2_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_2_cns_S0, shr_mem_2_cns_R0, shr_mem_2_cns_S1, shr_mem_2_cns_R1, shr_mem_2_cns_addra_shi0,
      shr_mem_2_cns_addra_shi1, shr_mem_2_cns_addrb_shi0, shr_mem_2_cns_addrb_shi1,
      shr_mem_2_cns_csa_n_shi0, shr_mem_2_cns_csa_n_shi1, shr_mem_2_cns_csb_n_shi0,
      shr_mem_2_cns_csb_n_shi1, shr_mem_2_cns_dinb_shi0, shr_mem_2_cns_dinb_shi1,
      shr_mem_2_cns_douta_sho0, shr_mem_2_cns_douta_sho1, shr_mem_2_cns_S1_pff, din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_2_cns_S0_pff
);
  input clk;
  input rst;
  input dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_2_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_2_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_2_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_2_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_2_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_2_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_2_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_2_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_2_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_2_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_2_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_2_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_2_cns_S0;
  input shr_mem_2_cns_R0;
  output shr_mem_2_cns_S1;
  input shr_mem_2_cns_R1;
  output [6:0] shr_mem_2_cns_addra_shi0;
  output [6:0] shr_mem_2_cns_addra_shi1;
  output [6:0] shr_mem_2_cns_addrb_shi0;
  output [6:0] shr_mem_2_cns_addrb_shi1;
  output shr_mem_2_cns_csa_n_shi0;
  output shr_mem_2_cns_csa_n_shi1;
  output shr_mem_2_cns_csb_n_shi0;
  output shr_mem_2_cns_csb_n_shi1;
  output [63:0] shr_mem_2_cns_dinb_shi0;
  output [63:0] shr_mem_2_cns_dinb_shi1;
  input [63:0] shr_mem_2_cns_douta_sho0;
  input [63:0] shr_mem_2_cns_douta_sho1;
  output shr_mem_2_cns_S1_pff;
  input din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_2_cns_S0_pff;


  // Interconnect Declarations
  reg dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_2_cns_PC0;
  reg shr_mem_2_cns_ppidx;
  reg [1:0] shr_mem_2_cns_ppown;
  wire shr_mem_2_cns_PC1;
  reg shr_mem_2_cns_ppidx_1;
  reg [1:0] shr_mem_2_cns_ppown_1;
  wire [6:0] shr_mem_2_shr_mem_2_mux_3_cse_pff;
  wire shr_mem_2_and_3_cse_pff;
  wire [1:0] shr_mem_2_acc_1_rmff;
  wire [3:0] nl_shr_mem_2_acc_1_rmff;
  wire shr_mem_2_xor_1_rmff;
  wire shr_mem_2_shr_mem_2_or_cse_pff;
  wire [1:0] shr_mem_2_acc_rmff;
  wire [3:0] nl_shr_mem_2_acc_rmff;
  wire shr_mem_2_xor_rmff;
  wire [6:0] shr_mem_2_shr_mem_2_mux_2_cse_pff;
  wire shr_mem_2_and_5_cse_pff;
  wire shr_mem_2_shr_mem_2_or_1_cse_pff;

  wire[0:0] shr_mem_2_mux_6_nl;
  wire[0:0] shr_mem_2_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_2_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_2_cns_R0;
  assign din_2_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_2_cns_R1;
  assign shr_mem_2_xor_rmff = shr_mem_2_cns_ppidx ^ shr_mem_2_cns_PC0;
  assign nl_shr_mem_2_acc_rmff = shr_mem_2_cns_ppown + conv_u2u_1_2(shr_mem_2_cns_PC0)
      + conv_s2u_1_2(shr_mem_2_cns_PC1);
  assign shr_mem_2_acc_rmff = nl_shr_mem_2_acc_rmff[1:0];
  assign shr_mem_2_cns_PC0 = shr_mem_2_cns_S0 & dout_2_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_2_xor_1_rmff = shr_mem_2_cns_ppidx_1 ^ shr_mem_2_cns_PC1;
  assign nl_shr_mem_2_acc_1_rmff = shr_mem_2_cns_ppown_1 + conv_u2u_1_2(shr_mem_2_cns_PC1)
      + conv_s2u_1_2(shr_mem_2_cns_PC0);
  assign shr_mem_2_acc_1_rmff = nl_shr_mem_2_acc_1_rmff[1:0];
  assign shr_mem_2_cns_PC1 = shr_mem_2_cns_S1 & din_2_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_2_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_2_cns_douta_sho0,
      shr_mem_2_cns_douta_sho1, shr_mem_2_cns_ppidx);
  assign din_2_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_2_cns_douta_sho0,
      shr_mem_2_cns_douta_sho1, shr_mem_2_cns_ppidx_1);
  assign shr_mem_2_cns_addra_shi0 = shr_mem_2_shr_mem_2_mux_3_cse_pff;
  assign shr_mem_2_cns_S1 = (shr_mem_2_cns_ppown_1!=2'b00);
  assign shr_mem_2_cns_S1_pff = (shr_mem_2_acc_1_rmff!=2'b00);
  assign shr_mem_2_and_3_cse_pff = shr_mem_2_cns_S1_pff & (~ shr_mem_2_xor_1_rmff);
  assign shr_mem_2_shr_mem_2_mux_3_cse_pff = MUX_v_7_2_2(dout_2_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_2_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_2_and_3_cse_pff);
  assign shr_mem_2_cns_addrb_shi0 = shr_mem_2_shr_mem_2_mux_3_cse_pff;
  assign shr_mem_2_cns_csa_n_shi0 = shr_mem_2_shr_mem_2_or_cse_pff;
  assign din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff = din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff = dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_2_cns_S0 = ~((shr_mem_2_cns_ppown==2'b10));
  assign shr_mem_2_cns_S0_pff = ~((shr_mem_2_acc_rmff==2'b10));
  assign shr_mem_2_mux_6_nl = MUX_s_1_2_2(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_2_and_3_cse_pff);
  assign shr_mem_2_shr_mem_2_or_cse_pff = (shr_mem_2_mux_6_nl) | (~((shr_mem_2_cns_S0_pff
      & (~ shr_mem_2_xor_rmff)) | shr_mem_2_and_3_cse_pff));
  assign shr_mem_2_cns_csb_n_shi0 = shr_mem_2_shr_mem_2_or_cse_pff;
  assign shr_mem_2_cns_dinb_shi0 = MUX_v_64_2_2(dout_2_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_2_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_2_and_3_cse_pff);
  assign shr_mem_2_cns_addra_shi1 = shr_mem_2_shr_mem_2_mux_2_cse_pff;
  assign shr_mem_2_and_5_cse_pff = shr_mem_2_cns_S1_pff & shr_mem_2_xor_1_rmff;
  assign shr_mem_2_shr_mem_2_mux_2_cse_pff = MUX_v_7_2_2(dout_2_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_2_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_2_and_5_cse_pff);
  assign shr_mem_2_cns_addrb_shi1 = shr_mem_2_shr_mem_2_mux_2_cse_pff;
  assign shr_mem_2_cns_csa_n_shi1 = shr_mem_2_shr_mem_2_or_1_cse_pff;
  assign shr_mem_2_mux_7_nl = MUX_s_1_2_2(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_2_and_5_cse_pff);
  assign shr_mem_2_shr_mem_2_or_1_cse_pff = (shr_mem_2_mux_7_nl) | (~((shr_mem_2_cns_S0_pff
      & shr_mem_2_xor_rmff) | shr_mem_2_and_5_cse_pff));
  assign shr_mem_2_cns_csb_n_shi1 = shr_mem_2_shr_mem_2_or_1_cse_pff;
  assign shr_mem_2_cns_dinb_shi1 = MUX_v_64_2_2(dout_2_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_2_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_2_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_2_cns_ppidx <= 1'b0;
      shr_mem_2_cns_ppown <= 2'b0;
      shr_mem_2_cns_ppidx_1 <= 1'b0;
      shr_mem_2_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_2_cns_ppidx <= shr_mem_2_xor_rmff;
      shr_mem_2_cns_ppown <= shr_mem_2_acc_rmff;
      shr_mem_2_cns_ppidx_1 <= shr_mem_2_xor_1_rmff;
      shr_mem_2_cns_ppown_1 <= shr_mem_2_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeaIgYu_1_cns_bctl
// ------------------------------------------------------------------


module double_buffeaIgYu_1_cns_bctl (
  clk, rst, dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_1_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_1_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_1_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_1_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_1_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_1_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_1_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_1_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_1_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_1_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_1_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_1_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_1_cns_S0, shr_mem_1_cns_R0, shr_mem_1_cns_S1, shr_mem_1_cns_R1, shr_mem_1_cns_addra_shi0,
      shr_mem_1_cns_addra_shi1, shr_mem_1_cns_addrb_shi0, shr_mem_1_cns_addrb_shi1,
      shr_mem_1_cns_csa_n_shi0, shr_mem_1_cns_csa_n_shi1, shr_mem_1_cns_csb_n_shi0,
      shr_mem_1_cns_csb_n_shi1, shr_mem_1_cns_dinb_shi0, shr_mem_1_cns_dinb_shi1,
      shr_mem_1_cns_douta_sho0, shr_mem_1_cns_douta_sho1, shr_mem_1_cns_S1_pff, din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff,
      din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff, dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff, shr_mem_1_cns_S0_pff
);
  input clk;
  input rst;
  input dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_1_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_1_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_1_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_1_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_1_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_1_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_1_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_1_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_1_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_1_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  output dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_1_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  output din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  output din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_1_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_1_cns_S0;
  input shr_mem_1_cns_R0;
  output shr_mem_1_cns_S1;
  input shr_mem_1_cns_R1;
  output [6:0] shr_mem_1_cns_addra_shi0;
  output [6:0] shr_mem_1_cns_addra_shi1;
  output [6:0] shr_mem_1_cns_addrb_shi0;
  output [6:0] shr_mem_1_cns_addrb_shi1;
  output shr_mem_1_cns_csa_n_shi0;
  output shr_mem_1_cns_csa_n_shi1;
  output shr_mem_1_cns_csb_n_shi0;
  output shr_mem_1_cns_csb_n_shi1;
  output [63:0] shr_mem_1_cns_dinb_shi0;
  output [63:0] shr_mem_1_cns_dinb_shi1;
  input [63:0] shr_mem_1_cns_douta_sho0;
  input [63:0] shr_mem_1_cns_douta_sho1;
  output shr_mem_1_cns_S1_pff;
  input din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  output din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  input dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  output dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output shr_mem_1_cns_S0_pff;


  // Interconnect Declarations
  reg dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  reg din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  reg din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  wire shr_mem_1_cns_PC0;
  reg shr_mem_1_cns_ppidx;
  reg [1:0] shr_mem_1_cns_ppown;
  wire shr_mem_1_cns_PC1;
  reg shr_mem_1_cns_ppidx_1;
  reg [1:0] shr_mem_1_cns_ppown_1;
  wire [6:0] shr_mem_1_shr_mem_1_mux_3_cse_pff;
  wire shr_mem_1_and_3_cse_pff;
  wire [1:0] shr_mem_1_acc_1_rmff;
  wire [3:0] nl_shr_mem_1_acc_1_rmff;
  wire shr_mem_1_xor_1_rmff;
  wire shr_mem_1_shr_mem_1_or_cse_pff;
  wire [1:0] shr_mem_1_acc_rmff;
  wire [3:0] nl_shr_mem_1_acc_rmff;
  wire shr_mem_1_xor_rmff;
  wire [6:0] shr_mem_1_shr_mem_1_mux_2_cse_pff;
  wire shr_mem_1_and_5_cse_pff;
  wire shr_mem_1_shr_mem_1_or_1_cse_pff;

  wire[0:0] shr_mem_1_mux_6_nl;
  wire[0:0] shr_mem_1_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign dout_1_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_1_cns_R0;
  assign din_1_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_1_cns_R1;
  assign shr_mem_1_xor_rmff = shr_mem_1_cns_ppidx ^ shr_mem_1_cns_PC0;
  assign nl_shr_mem_1_acc_rmff = shr_mem_1_cns_ppown + conv_u2u_1_2(shr_mem_1_cns_PC0)
      + conv_s2u_1_2(shr_mem_1_cns_PC1);
  assign shr_mem_1_acc_rmff = nl_shr_mem_1_acc_rmff[1:0];
  assign shr_mem_1_cns_PC0 = shr_mem_1_cns_S0 & dout_1_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_1_xor_1_rmff = shr_mem_1_cns_ppidx_1 ^ shr_mem_1_cns_PC1;
  assign nl_shr_mem_1_acc_1_rmff = shr_mem_1_cns_ppown_1 + conv_u2u_1_2(shr_mem_1_cns_PC1)
      + conv_s2u_1_2(shr_mem_1_cns_PC0);
  assign shr_mem_1_acc_1_rmff = nl_shr_mem_1_acc_1_rmff[1:0];
  assign shr_mem_1_cns_PC1 = shr_mem_1_cns_S1 & din_1_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_1_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_1_cns_douta_sho0,
      shr_mem_1_cns_douta_sho1, shr_mem_1_cns_ppidx);
  assign din_1_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_1_cns_douta_sho0,
      shr_mem_1_cns_douta_sho1, shr_mem_1_cns_ppidx_1);
  assign shr_mem_1_cns_addra_shi0 = shr_mem_1_shr_mem_1_mux_3_cse_pff;
  assign shr_mem_1_cns_S1 = (shr_mem_1_cns_ppown_1!=2'b00);
  assign shr_mem_1_cns_S1_pff = (shr_mem_1_acc_1_rmff!=2'b00);
  assign shr_mem_1_and_3_cse_pff = shr_mem_1_cns_S1_pff & (~ shr_mem_1_xor_1_rmff);
  assign shr_mem_1_shr_mem_1_mux_3_cse_pff = MUX_v_7_2_2(dout_1_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_1_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_1_and_3_cse_pff);
  assign shr_mem_1_cns_addrb_shi0 = shr_mem_1_shr_mem_1_mux_3_cse_pff;
  assign shr_mem_1_cns_csa_n_shi0 = shr_mem_1_shr_mem_1_or_cse_pff;
  assign din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud = ~ din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy;
  assign din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff = din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud = ~ dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy;
  assign dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff = dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign shr_mem_1_cns_S0 = ~((shr_mem_1_cns_ppown==2'b10));
  assign shr_mem_1_cns_S0_pff = ~((shr_mem_1_acc_rmff==2'b10));
  assign shr_mem_1_mux_6_nl = MUX_s_1_2_2(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_1_and_3_cse_pff);
  assign shr_mem_1_shr_mem_1_or_cse_pff = (shr_mem_1_mux_6_nl) | (~((shr_mem_1_cns_S0_pff
      & (~ shr_mem_1_xor_rmff)) | shr_mem_1_and_3_cse_pff));
  assign shr_mem_1_cns_csb_n_shi0 = shr_mem_1_shr_mem_1_or_cse_pff;
  assign shr_mem_1_cns_dinb_shi0 = MUX_v_64_2_2(dout_1_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_1_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_1_and_3_cse_pff);
  assign shr_mem_1_cns_addra_shi1 = shr_mem_1_shr_mem_1_mux_2_cse_pff;
  assign shr_mem_1_and_5_cse_pff = shr_mem_1_cns_S1_pff & shr_mem_1_xor_1_rmff;
  assign shr_mem_1_shr_mem_1_mux_2_cse_pff = MUX_v_7_2_2(dout_1_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_1_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_1_and_5_cse_pff);
  assign shr_mem_1_cns_addrb_shi1 = shr_mem_1_shr_mem_1_mux_2_cse_pff;
  assign shr_mem_1_cns_csa_n_shi1 = shr_mem_1_shr_mem_1_or_1_cse_pff;
  assign shr_mem_1_mux_7_nl = MUX_s_1_2_2(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff,
      din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, shr_mem_1_and_5_cse_pff);
  assign shr_mem_1_shr_mem_1_or_1_cse_pff = (shr_mem_1_mux_7_nl) | (~((shr_mem_1_cns_S0_pff
      & shr_mem_1_xor_rmff) | shr_mem_1_and_5_cse_pff));
  assign shr_mem_1_cns_csb_n_shi1 = shr_mem_1_shr_mem_1_or_1_cse_pff;
  assign shr_mem_1_cns_dinb_shi1 = MUX_v_64_2_2(dout_1_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_1_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_1_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= 1'b0;
      din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= 1'b0;
      shr_mem_1_cns_ppidx <= 1'b0;
      shr_mem_1_cns_ppown <= 2'b0;
      shr_mem_1_cns_ppidx_1 <= 1'b0;
      shr_mem_1_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buy <= ~ dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
      din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buy <= ~ din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
      shr_mem_1_cns_ppidx <= shr_mem_1_xor_rmff;
      shr_mem_1_cns_ppown <= shr_mem_1_acc_rmff;
      shr_mem_1_cns_ppidx_1 <= shr_mem_1_xor_1_rmff;
      shr_mem_1_cns_ppown_1 <= shr_mem_1_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeaIgYu_0_cns_bctl
// ------------------------------------------------------------------


module double_buffeaIgYu_0_cns_bctl (
  clk, rst, din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_0_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_0_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_0_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_0_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_0_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_0_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst, dout_0_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz, dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz, dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz, dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz, dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz, dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz, dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz, dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz, dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz,
      dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz, din_0_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_0_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_0_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_0_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_0_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      din_0_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_0_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst,
      dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz, din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz, din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz, din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz, din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz, din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz, din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz, din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz, din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz,
      din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud, dout_0_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_0_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_1_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_1_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_2_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_2_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_3_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_3_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_4_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_4_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_5_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_5_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_6_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_6_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_7_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_7_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_8_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_8_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_9_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_9_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_10_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_10_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_11_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_11_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_12_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_12_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_13_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_13_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_14_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_14_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_15_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_15_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_16_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_16_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud,
      dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud, dout_17_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud,
      din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud, din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud,
      din_17_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud, dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud,
      shr_mem_0_cns_S0, shr_mem_0_cns_R0, shr_mem_0_cns_S1, shr_mem_0_cns_R1, shr_mem_0_cns_addra_shi0,
      shr_mem_0_cns_addra_shi1, shr_mem_0_cns_addrb_shi0, shr_mem_0_cns_addrb_shi1,
      shr_mem_0_cns_csa_n_shi0, shr_mem_0_cns_csa_n_shi1, shr_mem_0_cns_csb_n_shi0,
      shr_mem_0_cns_csb_n_shi1, shr_mem_0_cns_dinb_shi0, shr_mem_0_cns_dinb_shi1,
      shr_mem_0_cns_douta_sho0, shr_mem_0_cns_douta_sho1, shr_mem_0_cns_S1_pff, shr_mem_0_cns_S0_pff,
      din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff,
      din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff, din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff,
      dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff, dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff
);
  input clk;
  input rst;
  output din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_0_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input dout_0_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_0_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [6:0] dout_0_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  input [63:0] dout_0_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output [63:0] dout_0_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_0_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  output dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  output dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  input din_0_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input din_0_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_0_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [6:0] din_0_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  input [63:0] din_0_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output [63:0] din_0_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_0_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  output din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  output din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  input din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input dout_0_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_0_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_1_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_1_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_2_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_2_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_3_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_3_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_4_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_4_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_5_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_5_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_6_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_6_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_7_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_7_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_8_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_8_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_9_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_9_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_10_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_10_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_11_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_11_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_12_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_12_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_13_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_13_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_14_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_14_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_15_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_15_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_16_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_16_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  input dout_17_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  input din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  input din_17_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  input dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  output shr_mem_0_cns_S0;
  input shr_mem_0_cns_R0;
  output shr_mem_0_cns_S1;
  input shr_mem_0_cns_R1;
  output [6:0] shr_mem_0_cns_addra_shi0;
  output [6:0] shr_mem_0_cns_addra_shi1;
  output [6:0] shr_mem_0_cns_addrb_shi0;
  output [6:0] shr_mem_0_cns_addrb_shi1;
  output shr_mem_0_cns_csa_n_shi0;
  output shr_mem_0_cns_csa_n_shi1;
  output shr_mem_0_cns_csb_n_shi0;
  output shr_mem_0_cns_csb_n_shi1;
  output [63:0] shr_mem_0_cns_dinb_shi0;
  output [63:0] shr_mem_0_cns_dinb_shi1;
  input [63:0] shr_mem_0_cns_douta_sho0;
  input [63:0] shr_mem_0_cns_douta_sho1;
  output shr_mem_0_cns_S1_pff;
  output shr_mem_0_cns_S0_pff;
  output din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  output din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff;
  input din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  output dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff;
  input dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;


  // Interconnect Declarations
  wire shr_mem_0_cns_PC0;
  reg shr_mem_0_cns_ppidx;
  reg [1:0] shr_mem_0_cns_ppown;
  wire shr_mem_0_cns_PC1;
  reg shr_mem_0_cns_ppidx_1;
  reg [1:0] shr_mem_0_cns_ppown_1;
  wire [6:0] shr_mem_0_shr_mem_0_mux_3_cse_pff;
  wire shr_mem_0_and_3_cse_pff;
  wire [1:0] shr_mem_0_acc_1_rmff;
  wire [3:0] nl_shr_mem_0_acc_1_rmff;
  wire shr_mem_0_xor_1_rmff;
  wire shr_mem_0_shr_mem_0_shr_mem_0_nand_cse_pff;
  wire [1:0] shr_mem_0_acc_rmff;
  wire [3:0] nl_shr_mem_0_acc_rmff;
  wire shr_mem_0_xor_rmff;
  wire [6:0] shr_mem_0_shr_mem_0_mux_2_cse_pff;
  wire shr_mem_0_and_5_cse_pff;
  wire shr_mem_0_shr_mem_0_shr_mem_0_nand_1_cse_pff;

  wire[0:0] shr_mem_0_mux_6_nl;
  wire[0:0] shr_mem_0_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_0_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = shr_mem_0_cns_R0;
  assign din_0_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = shr_mem_0_cns_R1;
  assign shr_mem_0_xor_rmff = shr_mem_0_cns_ppidx ^ shr_mem_0_cns_PC0;
  assign nl_shr_mem_0_acc_rmff = shr_mem_0_cns_ppown + conv_u2u_1_2(shr_mem_0_cns_PC0)
      + conv_s2u_1_2(shr_mem_0_cns_PC1);
  assign shr_mem_0_acc_rmff = nl_shr_mem_0_acc_rmff[1:0];
  assign shr_mem_0_cns_PC0 = shr_mem_0_cns_S0 & dout_0_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  assign shr_mem_0_xor_1_rmff = shr_mem_0_cns_ppidx_1 ^ shr_mem_0_cns_PC1;
  assign nl_shr_mem_0_acc_1_rmff = shr_mem_0_cns_ppown_1 + conv_u2u_1_2(shr_mem_0_cns_PC1)
      + conv_s2u_1_2(shr_mem_0_cns_PC0);
  assign shr_mem_0_acc_1_rmff = nl_shr_mem_0_acc_1_rmff[1:0];
  assign shr_mem_0_cns_PC1 = shr_mem_0_cns_S1 & din_0_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  assign dout_0_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst = MUX_v_64_2_2(shr_mem_0_cns_douta_sho0,
      shr_mem_0_cns_douta_sho1, shr_mem_0_cns_ppidx);
  assign din_0_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst = MUX_v_64_2_2(shr_mem_0_cns_douta_sho0,
      shr_mem_0_cns_douta_sho1, shr_mem_0_cns_ppidx_1);
  assign shr_mem_0_cns_addra_shi0 = shr_mem_0_shr_mem_0_mux_3_cse_pff;
  assign shr_mem_0_cns_S1 = (shr_mem_0_cns_ppown_1!=2'b00);
  assign shr_mem_0_cns_S1_pff = (shr_mem_0_acc_1_rmff!=2'b00);
  assign shr_mem_0_and_3_cse_pff = shr_mem_0_cns_S1_pff & (~ shr_mem_0_xor_1_rmff);
  assign shr_mem_0_shr_mem_0_mux_3_cse_pff = MUX_v_7_2_2(dout_0_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_0_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_0_and_3_cse_pff);
  assign shr_mem_0_cns_addrb_shi0 = shr_mem_0_shr_mem_0_mux_3_cse_pff;
  assign shr_mem_0_cns_csa_n_shi0 = shr_mem_0_shr_mem_0_shr_mem_0_nand_cse_pff;
  assign shr_mem_0_cns_S0 = ~((shr_mem_0_cns_ppown==2'b10));
  assign shr_mem_0_cns_S0_pff = ~((shr_mem_0_acc_rmff==2'b10));
  assign shr_mem_0_mux_6_nl = MUX_s_1_2_2(dout_0_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_0_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_0_and_3_cse_pff);
  assign shr_mem_0_shr_mem_0_shr_mem_0_nand_cse_pff = (shr_mem_0_mux_6_nl) | (~((shr_mem_0_cns_S0_pff
      & (~ shr_mem_0_xor_rmff)) | shr_mem_0_and_3_cse_pff));
  assign shr_mem_0_cns_csb_n_shi0 = shr_mem_0_shr_mem_0_shr_mem_0_nand_cse_pff;
  assign shr_mem_0_cns_dinb_shi0 = MUX_v_64_2_2(dout_0_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_0_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_0_and_3_cse_pff);
  assign shr_mem_0_cns_addra_shi1 = shr_mem_0_shr_mem_0_mux_2_cse_pff;
  assign shr_mem_0_and_5_cse_pff = shr_mem_0_cns_S1_pff & shr_mem_0_xor_1_rmff;
  assign shr_mem_0_shr_mem_0_mux_2_cse_pff = MUX_v_7_2_2(dout_0_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_0_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_0_and_5_cse_pff);
  assign shr_mem_0_cns_addrb_shi1 = shr_mem_0_shr_mem_0_mux_2_cse_pff;
  assign shr_mem_0_cns_csa_n_shi1 = shr_mem_0_shr_mem_0_shr_mem_0_nand_1_cse_pff;
  assign shr_mem_0_mux_7_nl = MUX_s_1_2_2(dout_0_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_0_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_0_and_5_cse_pff);
  assign shr_mem_0_shr_mem_0_shr_mem_0_nand_1_cse_pff = (shr_mem_0_mux_7_nl) | (~((shr_mem_0_cns_S0_pff
      & shr_mem_0_xor_rmff) | shr_mem_0_and_5_cse_pff));
  assign shr_mem_0_cns_csb_n_shi1 = shr_mem_0_shr_mem_0_shr_mem_0_nand_1_cse_pff;
  assign shr_mem_0_cns_dinb_shi1 = MUX_v_64_2_2(dout_0_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst,
      din_0_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst, shr_mem_0_and_5_cse_pff);
  assign din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  assign din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz = din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  assign din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff = din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff;
  assign dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz = dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  assign dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff = dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff;
  always @(posedge clk) begin
    if ( rst ) begin
      shr_mem_0_cns_ppidx <= 1'b0;
      shr_mem_0_cns_ppown <= 2'b0;
      shr_mem_0_cns_ppidx_1 <= 1'b0;
      shr_mem_0_cns_ppown_1 <= 2'b0;
    end
    else begin
      shr_mem_0_cns_ppidx <= shr_mem_0_xor_rmff;
      shr_mem_0_cns_ppown <= shr_mem_0_acc_rmff;
      shr_mem_0_cns_ppidx_1 <= shr_mem_0_xor_1_rmff;
      shr_mem_0_cns_ppown_1 <= shr_mem_0_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    unreg_hier_69
// ------------------------------------------------------------------


module unreg_hier_69 (
  in_0, out_0
);
  input in_0;
  output out_0;



  // Interconnect Declarations for Component Instantiations 
  assign out_0 = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_37_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_37_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_17_data_and_nl;
  wire tmp_17_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_17_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_17_data_and_nl);
  assign tmp_17_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_17_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_36_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_36_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_16_data_and_nl;
  wire tmp_16_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_16_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_16_data_and_nl);
  assign tmp_16_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_16_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_35_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_35_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_15_data_and_nl;
  wire tmp_15_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_15_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_15_data_and_nl);
  assign tmp_15_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_15_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_34_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_34_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_14_data_and_nl;
  wire tmp_14_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_14_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_14_data_and_nl);
  assign tmp_14_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_14_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_33_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_33_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_13_data_and_nl;
  wire tmp_13_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_13_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_13_data_and_nl);
  assign tmp_13_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_13_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_32_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_32_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_12_data_and_nl;
  wire tmp_12_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_12_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_12_data_and_nl);
  assign tmp_12_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_12_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_31_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_31_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_11_data_and_nl;
  wire tmp_11_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_11_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_11_data_and_nl);
  assign tmp_11_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_11_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_30_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_30_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_10_data_and_nl;
  wire tmp_10_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_10_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_10_data_and_nl);
  assign tmp_10_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_10_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_29_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_29_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_9_data_and_nl;
  wire tmp_9_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_9_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_9_data_and_nl);
  assign tmp_9_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_9_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_28_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_28_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_8_data_and_nl;
  wire tmp_8_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_8_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_8_data_and_nl);
  assign tmp_8_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_8_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_27_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_27_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_7_data_and_nl;
  wire tmp_7_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_7_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_7_data_and_nl);
  assign tmp_7_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_7_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_26_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_26_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_6_data_and_nl;
  wire tmp_6_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_6_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_6_data_and_nl);
  assign tmp_6_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_6_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_25_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_25_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_5_data_and_nl;
  wire tmp_5_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_5_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_5_data_and_nl);
  assign tmp_5_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_5_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_24_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_24_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_4_data_and_nl;
  wire tmp_4_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_4_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_4_data_and_nl);
  assign tmp_4_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_4_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_23_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_23_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_3_data_and_nl;
  wire tmp_3_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_3_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_3_data_and_nl);
  assign tmp_3_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_3_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_22_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_22_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_2_data_and_nl;
  wire tmp_2_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_2_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_2_data_and_nl);
  assign tmp_2_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_2_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_21_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_21_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_1_data_and_nl;
  wire tmp_1_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_1_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_1_data_and_nl);
  assign tmp_1_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_1_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_20_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_20_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire tmp_0_data_and_nl;
  wire tmp_0_data_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign tmp_0_data_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (tmp_0_data_and_nl);
  assign tmp_0_data_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (tmp_0_data_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_19_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_19_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_17_and_nl;
  wire dout_17_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_17_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_17_and_nl);
  assign dout_17_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_17_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_18_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_18_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_16_and_nl;
  wire dout_16_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_16_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_16_and_nl);
  assign dout_16_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_16_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_17_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_17_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_15_and_nl;
  wire dout_15_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_15_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_15_and_nl);
  assign dout_15_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_15_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_16_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_16_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_14_and_nl;
  wire dout_14_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_14_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_14_and_nl);
  assign dout_14_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_14_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_15_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_15_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_13_and_nl;
  wire dout_13_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_13_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_13_and_nl);
  assign dout_13_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_13_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_14_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_14_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_12_and_nl;
  wire dout_12_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_12_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_12_and_nl);
  assign dout_12_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_12_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_13_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_13_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_11_and_nl;
  wire dout_11_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_11_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_11_and_nl);
  assign dout_11_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_11_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_12_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_12_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_10_and_nl;
  wire dout_10_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_10_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_10_and_nl);
  assign dout_10_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_10_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_11_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_11_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_9_and_nl;
  wire dout_9_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_9_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_9_and_nl);
  assign dout_9_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_9_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_10_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_10_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_8_and_nl;
  wire dout_8_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_8_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_8_and_nl);
  assign dout_8_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_8_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_9_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_9_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_7_and_nl;
  wire dout_7_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_7_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_7_and_nl);
  assign dout_7_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_7_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_8_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_8_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_6_and_nl;
  wire dout_6_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_6_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_6_and_nl);
  assign dout_6_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_6_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_7_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_7_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_5_and_nl;
  wire dout_5_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_5_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_5_and_nl);
  assign dout_5_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_5_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_6_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_6_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_4_and_nl;
  wire dout_4_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_4_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_4_and_nl);
  assign dout_4_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_4_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_5_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_5_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_3_and_nl;
  wire dout_3_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_3_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_3_and_nl);
  assign dout_3_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_3_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_4_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_4_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_2_and_nl;
  wire dout_2_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_2_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_2_and_nl);
  assign dout_2_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_2_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_3_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_3_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_1_and_nl;
  wire dout_1_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_1_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_1_and_nl);
  assign dout_1_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_1_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_2_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_2_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_0_and_nl;
  wire dout_0_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_0_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_0_and_nl);
  assign dout_0_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_0_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_staller
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_staller (
  clk, rst, core_wen, din_rsci_wen_comp, core_wten, dout_17_rsc_req_obj_wen_comp,
      dout_16_rsc_req_obj_wen_comp, dout_15_rsc_req_obj_wen_comp, dout_14_rsc_req_obj_wen_comp,
      dout_13_rsc_req_obj_wen_comp, dout_12_rsc_req_obj_wen_comp, dout_11_rsc_req_obj_wen_comp,
      dout_10_rsc_req_obj_wen_comp, dout_9_rsc_req_obj_wen_comp, dout_8_rsc_req_obj_wen_comp,
      dout_7_rsc_req_obj_wen_comp, dout_6_rsc_req_obj_wen_comp, dout_5_rsc_req_obj_wen_comp,
      dout_4_rsc_req_obj_wen_comp, dout_3_rsc_req_obj_wen_comp, dout_2_rsc_req_obj_wen_comp,
      dout_1_rsc_req_obj_wen_comp, dout_0_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  input din_rsci_wen_comp;
  output core_wten;
  input dout_17_rsc_req_obj_wen_comp;
  input dout_16_rsc_req_obj_wen_comp;
  input dout_15_rsc_req_obj_wen_comp;
  input dout_14_rsc_req_obj_wen_comp;
  input dout_13_rsc_req_obj_wen_comp;
  input dout_12_rsc_req_obj_wen_comp;
  input dout_11_rsc_req_obj_wen_comp;
  input dout_10_rsc_req_obj_wen_comp;
  input dout_9_rsc_req_obj_wen_comp;
  input dout_8_rsc_req_obj_wen_comp;
  input dout_7_rsc_req_obj_wen_comp;
  input dout_6_rsc_req_obj_wen_comp;
  input dout_5_rsc_req_obj_wen_comp;
  input dout_4_rsc_req_obj_wen_comp;
  input dout_3_rsc_req_obj_wen_comp;
  input dout_2_rsc_req_obj_wen_comp;
  input dout_1_rsc_req_obj_wen_comp;
  input dout_0_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = din_rsci_wen_comp & dout_17_rsc_req_obj_wen_comp & dout_16_rsc_req_obj_wen_comp
      & dout_15_rsc_req_obj_wen_comp & dout_14_rsc_req_obj_wen_comp & dout_13_rsc_req_obj_wen_comp
      & dout_12_rsc_req_obj_wen_comp & dout_11_rsc_req_obj_wen_comp & dout_10_rsc_req_obj_wen_comp
      & dout_9_rsc_req_obj_wen_comp & dout_8_rsc_req_obj_wen_comp & dout_7_rsc_req_obj_wen_comp
      & dout_6_rsc_req_obj_wen_comp & dout_5_rsc_req_obj_wen_comp & dout_4_rsc_req_obj_wen_comp
      & dout_3_rsc_req_obj_wen_comp & dout_2_rsc_req_obj_wen_comp & dout_1_rsc_req_obj_wen_comp
      & dout_0_rsc_req_obj_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_dp
    (
  clk, rst, dout_0_rsc_req_obj_oswt, dout_0_rsc_req_obj_wen_comp, dout_0_rsc_req_obj_biwt,
      dout_0_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_0_rsc_req_obj_oswt;
  output dout_0_rsc_req_obj_wen_comp;
  input dout_0_rsc_req_obj_biwt;
  input dout_0_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_0_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_0_rsc_req_obj_wen_comp = (~ dout_0_rsc_req_obj_oswt) | dout_0_rsc_req_obj_biwt
      | dout_0_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_0_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_0_rsc_req_obj_bcwt <= ~((~(dout_0_rsc_req_obj_bcwt | dout_0_rsc_req_obj_biwt))
          | dout_0_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_0_rsc_req_obj_oswt, dout_0_rsc_req_obj_vd,
      dout_0_rsc_req_obj_biwt, dout_0_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_0_rsc_req_obj_oswt;
  input dout_0_rsc_req_obj_vd;
  output dout_0_rsc_req_obj_biwt;
  output dout_0_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_0_rsc_req_obj_pdswt0;
  reg dout_0_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_0_rsc_req_obj_pdswt0 = (~ core_wten) & dout_0_rsc_req_obj_oswt;
  assign dout_0_rsc_req_obj_biwt = (dout_0_rsc_req_obj_pdswt0 | dout_0_rsc_req_obj_icwt)
      & dout_0_rsc_req_obj_vd;
  assign dout_0_rsc_req_obj_bdwt = dout_0_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_0_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_0_rsc_req_obj_icwt <= ~((~(dout_0_rsc_req_obj_icwt | dout_0_rsc_req_obj_pdswt0))
          | dout_0_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_rls_obj_dout_0_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_rls_obj_dout_0_rsc_rls_wait_ctrl
    (
  core_wten, dout_0_rsc_rls_obj_iswt0, dout_0_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_0_rsc_rls_obj_iswt0;
  output dout_0_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_0_rsc_rls_obj_ld_core_sct = dout_0_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_dp
    (
  clk, rst, dout_1_rsc_req_obj_oswt, dout_1_rsc_req_obj_wen_comp, dout_1_rsc_req_obj_biwt,
      dout_1_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_1_rsc_req_obj_oswt;
  output dout_1_rsc_req_obj_wen_comp;
  input dout_1_rsc_req_obj_biwt;
  input dout_1_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_1_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_1_rsc_req_obj_wen_comp = (~ dout_1_rsc_req_obj_oswt) | dout_1_rsc_req_obj_biwt
      | dout_1_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_1_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_1_rsc_req_obj_bcwt <= ~((~(dout_1_rsc_req_obj_bcwt | dout_1_rsc_req_obj_biwt))
          | dout_1_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_1_rsc_req_obj_oswt, dout_1_rsc_req_obj_vd,
      dout_1_rsc_req_obj_biwt, dout_1_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_1_rsc_req_obj_oswt;
  input dout_1_rsc_req_obj_vd;
  output dout_1_rsc_req_obj_biwt;
  output dout_1_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_1_rsc_req_obj_pdswt0;
  reg dout_1_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_1_rsc_req_obj_pdswt0 = (~ core_wten) & dout_1_rsc_req_obj_oswt;
  assign dout_1_rsc_req_obj_biwt = (dout_1_rsc_req_obj_pdswt0 | dout_1_rsc_req_obj_icwt)
      & dout_1_rsc_req_obj_vd;
  assign dout_1_rsc_req_obj_bdwt = dout_1_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_1_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_1_rsc_req_obj_icwt <= ~((~(dout_1_rsc_req_obj_icwt | dout_1_rsc_req_obj_pdswt0))
          | dout_1_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_rls_obj_dout_1_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_rls_obj_dout_1_rsc_rls_wait_ctrl
    (
  core_wten, dout_1_rsc_rls_obj_iswt0, dout_1_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_1_rsc_rls_obj_iswt0;
  output dout_1_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_1_rsc_rls_obj_ld_core_sct = dout_1_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_dp
    (
  clk, rst, dout_2_rsc_req_obj_oswt, dout_2_rsc_req_obj_wen_comp, dout_2_rsc_req_obj_biwt,
      dout_2_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_2_rsc_req_obj_oswt;
  output dout_2_rsc_req_obj_wen_comp;
  input dout_2_rsc_req_obj_biwt;
  input dout_2_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_2_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_2_rsc_req_obj_wen_comp = (~ dout_2_rsc_req_obj_oswt) | dout_2_rsc_req_obj_biwt
      | dout_2_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_2_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_2_rsc_req_obj_bcwt <= ~((~(dout_2_rsc_req_obj_bcwt | dout_2_rsc_req_obj_biwt))
          | dout_2_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_2_rsc_req_obj_oswt, dout_2_rsc_req_obj_vd,
      dout_2_rsc_req_obj_biwt, dout_2_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_2_rsc_req_obj_oswt;
  input dout_2_rsc_req_obj_vd;
  output dout_2_rsc_req_obj_biwt;
  output dout_2_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_2_rsc_req_obj_pdswt0;
  reg dout_2_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_2_rsc_req_obj_pdswt0 = (~ core_wten) & dout_2_rsc_req_obj_oswt;
  assign dout_2_rsc_req_obj_biwt = (dout_2_rsc_req_obj_pdswt0 | dout_2_rsc_req_obj_icwt)
      & dout_2_rsc_req_obj_vd;
  assign dout_2_rsc_req_obj_bdwt = dout_2_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_2_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_2_rsc_req_obj_icwt <= ~((~(dout_2_rsc_req_obj_icwt | dout_2_rsc_req_obj_pdswt0))
          | dout_2_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_rls_obj_dout_2_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_rls_obj_dout_2_rsc_rls_wait_ctrl
    (
  core_wten, dout_2_rsc_rls_obj_iswt0, dout_2_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_2_rsc_rls_obj_iswt0;
  output dout_2_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_2_rsc_rls_obj_ld_core_sct = dout_2_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_dp
    (
  clk, rst, dout_3_rsc_req_obj_oswt, dout_3_rsc_req_obj_wen_comp, dout_3_rsc_req_obj_biwt,
      dout_3_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_3_rsc_req_obj_oswt;
  output dout_3_rsc_req_obj_wen_comp;
  input dout_3_rsc_req_obj_biwt;
  input dout_3_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_3_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_3_rsc_req_obj_wen_comp = (~ dout_3_rsc_req_obj_oswt) | dout_3_rsc_req_obj_biwt
      | dout_3_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_3_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_3_rsc_req_obj_bcwt <= ~((~(dout_3_rsc_req_obj_bcwt | dout_3_rsc_req_obj_biwt))
          | dout_3_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_3_rsc_req_obj_oswt, dout_3_rsc_req_obj_vd,
      dout_3_rsc_req_obj_biwt, dout_3_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_3_rsc_req_obj_oswt;
  input dout_3_rsc_req_obj_vd;
  output dout_3_rsc_req_obj_biwt;
  output dout_3_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_3_rsc_req_obj_pdswt0;
  reg dout_3_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_3_rsc_req_obj_pdswt0 = (~ core_wten) & dout_3_rsc_req_obj_oswt;
  assign dout_3_rsc_req_obj_biwt = (dout_3_rsc_req_obj_pdswt0 | dout_3_rsc_req_obj_icwt)
      & dout_3_rsc_req_obj_vd;
  assign dout_3_rsc_req_obj_bdwt = dout_3_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_3_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_3_rsc_req_obj_icwt <= ~((~(dout_3_rsc_req_obj_icwt | dout_3_rsc_req_obj_pdswt0))
          | dout_3_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_rls_obj_dout_3_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_rls_obj_dout_3_rsc_rls_wait_ctrl
    (
  core_wten, dout_3_rsc_rls_obj_iswt0, dout_3_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_3_rsc_rls_obj_iswt0;
  output dout_3_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_3_rsc_rls_obj_ld_core_sct = dout_3_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_dp
    (
  clk, rst, dout_4_rsc_req_obj_oswt, dout_4_rsc_req_obj_wen_comp, dout_4_rsc_req_obj_biwt,
      dout_4_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_4_rsc_req_obj_oswt;
  output dout_4_rsc_req_obj_wen_comp;
  input dout_4_rsc_req_obj_biwt;
  input dout_4_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_4_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_4_rsc_req_obj_wen_comp = (~ dout_4_rsc_req_obj_oswt) | dout_4_rsc_req_obj_biwt
      | dout_4_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_4_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_4_rsc_req_obj_bcwt <= ~((~(dout_4_rsc_req_obj_bcwt | dout_4_rsc_req_obj_biwt))
          | dout_4_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_4_rsc_req_obj_oswt, dout_4_rsc_req_obj_vd,
      dout_4_rsc_req_obj_biwt, dout_4_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_4_rsc_req_obj_oswt;
  input dout_4_rsc_req_obj_vd;
  output dout_4_rsc_req_obj_biwt;
  output dout_4_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_4_rsc_req_obj_pdswt0;
  reg dout_4_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_4_rsc_req_obj_pdswt0 = (~ core_wten) & dout_4_rsc_req_obj_oswt;
  assign dout_4_rsc_req_obj_biwt = (dout_4_rsc_req_obj_pdswt0 | dout_4_rsc_req_obj_icwt)
      & dout_4_rsc_req_obj_vd;
  assign dout_4_rsc_req_obj_bdwt = dout_4_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_4_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_4_rsc_req_obj_icwt <= ~((~(dout_4_rsc_req_obj_icwt | dout_4_rsc_req_obj_pdswt0))
          | dout_4_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_rls_obj_dout_4_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_rls_obj_dout_4_rsc_rls_wait_ctrl
    (
  core_wten, dout_4_rsc_rls_obj_iswt0, dout_4_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_4_rsc_rls_obj_iswt0;
  output dout_4_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_4_rsc_rls_obj_ld_core_sct = dout_4_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_dp
    (
  clk, rst, dout_5_rsc_req_obj_oswt, dout_5_rsc_req_obj_wen_comp, dout_5_rsc_req_obj_biwt,
      dout_5_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_5_rsc_req_obj_oswt;
  output dout_5_rsc_req_obj_wen_comp;
  input dout_5_rsc_req_obj_biwt;
  input dout_5_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_5_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_5_rsc_req_obj_wen_comp = (~ dout_5_rsc_req_obj_oswt) | dout_5_rsc_req_obj_biwt
      | dout_5_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_5_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_5_rsc_req_obj_bcwt <= ~((~(dout_5_rsc_req_obj_bcwt | dout_5_rsc_req_obj_biwt))
          | dout_5_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_5_rsc_req_obj_oswt, dout_5_rsc_req_obj_vd,
      dout_5_rsc_req_obj_biwt, dout_5_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_5_rsc_req_obj_oswt;
  input dout_5_rsc_req_obj_vd;
  output dout_5_rsc_req_obj_biwt;
  output dout_5_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_5_rsc_req_obj_pdswt0;
  reg dout_5_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_5_rsc_req_obj_pdswt0 = (~ core_wten) & dout_5_rsc_req_obj_oswt;
  assign dout_5_rsc_req_obj_biwt = (dout_5_rsc_req_obj_pdswt0 | dout_5_rsc_req_obj_icwt)
      & dout_5_rsc_req_obj_vd;
  assign dout_5_rsc_req_obj_bdwt = dout_5_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_5_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_5_rsc_req_obj_icwt <= ~((~(dout_5_rsc_req_obj_icwt | dout_5_rsc_req_obj_pdswt0))
          | dout_5_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_rls_obj_dout_5_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_rls_obj_dout_5_rsc_rls_wait_ctrl
    (
  core_wten, dout_5_rsc_rls_obj_iswt0, dout_5_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_5_rsc_rls_obj_iswt0;
  output dout_5_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_5_rsc_rls_obj_ld_core_sct = dout_5_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_dp
    (
  clk, rst, dout_6_rsc_req_obj_oswt, dout_6_rsc_req_obj_wen_comp, dout_6_rsc_req_obj_biwt,
      dout_6_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_6_rsc_req_obj_oswt;
  output dout_6_rsc_req_obj_wen_comp;
  input dout_6_rsc_req_obj_biwt;
  input dout_6_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_6_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_6_rsc_req_obj_wen_comp = (~ dout_6_rsc_req_obj_oswt) | dout_6_rsc_req_obj_biwt
      | dout_6_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_6_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_6_rsc_req_obj_bcwt <= ~((~(dout_6_rsc_req_obj_bcwt | dout_6_rsc_req_obj_biwt))
          | dout_6_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_6_rsc_req_obj_oswt, dout_6_rsc_req_obj_vd,
      dout_6_rsc_req_obj_biwt, dout_6_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_6_rsc_req_obj_oswt;
  input dout_6_rsc_req_obj_vd;
  output dout_6_rsc_req_obj_biwt;
  output dout_6_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_6_rsc_req_obj_pdswt0;
  reg dout_6_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_6_rsc_req_obj_pdswt0 = (~ core_wten) & dout_6_rsc_req_obj_oswt;
  assign dout_6_rsc_req_obj_biwt = (dout_6_rsc_req_obj_pdswt0 | dout_6_rsc_req_obj_icwt)
      & dout_6_rsc_req_obj_vd;
  assign dout_6_rsc_req_obj_bdwt = dout_6_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_6_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_6_rsc_req_obj_icwt <= ~((~(dout_6_rsc_req_obj_icwt | dout_6_rsc_req_obj_pdswt0))
          | dout_6_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_rls_obj_dout_6_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_rls_obj_dout_6_rsc_rls_wait_ctrl
    (
  core_wten, dout_6_rsc_rls_obj_iswt0, dout_6_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_6_rsc_rls_obj_iswt0;
  output dout_6_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_6_rsc_rls_obj_ld_core_sct = dout_6_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_dp
    (
  clk, rst, dout_7_rsc_req_obj_oswt, dout_7_rsc_req_obj_wen_comp, dout_7_rsc_req_obj_biwt,
      dout_7_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_7_rsc_req_obj_oswt;
  output dout_7_rsc_req_obj_wen_comp;
  input dout_7_rsc_req_obj_biwt;
  input dout_7_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_7_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_7_rsc_req_obj_wen_comp = (~ dout_7_rsc_req_obj_oswt) | dout_7_rsc_req_obj_biwt
      | dout_7_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_7_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_7_rsc_req_obj_bcwt <= ~((~(dout_7_rsc_req_obj_bcwt | dout_7_rsc_req_obj_biwt))
          | dout_7_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_7_rsc_req_obj_oswt, dout_7_rsc_req_obj_vd,
      dout_7_rsc_req_obj_biwt, dout_7_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_7_rsc_req_obj_oswt;
  input dout_7_rsc_req_obj_vd;
  output dout_7_rsc_req_obj_biwt;
  output dout_7_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_7_rsc_req_obj_pdswt0;
  reg dout_7_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_7_rsc_req_obj_pdswt0 = (~ core_wten) & dout_7_rsc_req_obj_oswt;
  assign dout_7_rsc_req_obj_biwt = (dout_7_rsc_req_obj_pdswt0 | dout_7_rsc_req_obj_icwt)
      & dout_7_rsc_req_obj_vd;
  assign dout_7_rsc_req_obj_bdwt = dout_7_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_7_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_7_rsc_req_obj_icwt <= ~((~(dout_7_rsc_req_obj_icwt | dout_7_rsc_req_obj_pdswt0))
          | dout_7_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_rls_obj_dout_7_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_rls_obj_dout_7_rsc_rls_wait_ctrl
    (
  core_wten, dout_7_rsc_rls_obj_iswt0, dout_7_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_7_rsc_rls_obj_iswt0;
  output dout_7_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_7_rsc_rls_obj_ld_core_sct = dout_7_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_dp
    (
  clk, rst, dout_8_rsc_req_obj_oswt, dout_8_rsc_req_obj_wen_comp, dout_8_rsc_req_obj_biwt,
      dout_8_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_8_rsc_req_obj_oswt;
  output dout_8_rsc_req_obj_wen_comp;
  input dout_8_rsc_req_obj_biwt;
  input dout_8_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_8_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_8_rsc_req_obj_wen_comp = (~ dout_8_rsc_req_obj_oswt) | dout_8_rsc_req_obj_biwt
      | dout_8_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_8_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_8_rsc_req_obj_bcwt <= ~((~(dout_8_rsc_req_obj_bcwt | dout_8_rsc_req_obj_biwt))
          | dout_8_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_8_rsc_req_obj_oswt, dout_8_rsc_req_obj_vd,
      dout_8_rsc_req_obj_biwt, dout_8_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_8_rsc_req_obj_oswt;
  input dout_8_rsc_req_obj_vd;
  output dout_8_rsc_req_obj_biwt;
  output dout_8_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_8_rsc_req_obj_pdswt0;
  reg dout_8_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_8_rsc_req_obj_pdswt0 = (~ core_wten) & dout_8_rsc_req_obj_oswt;
  assign dout_8_rsc_req_obj_biwt = (dout_8_rsc_req_obj_pdswt0 | dout_8_rsc_req_obj_icwt)
      & dout_8_rsc_req_obj_vd;
  assign dout_8_rsc_req_obj_bdwt = dout_8_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_8_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_8_rsc_req_obj_icwt <= ~((~(dout_8_rsc_req_obj_icwt | dout_8_rsc_req_obj_pdswt0))
          | dout_8_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_rls_obj_dout_8_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_rls_obj_dout_8_rsc_rls_wait_ctrl
    (
  core_wten, dout_8_rsc_rls_obj_iswt0, dout_8_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_8_rsc_rls_obj_iswt0;
  output dout_8_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_8_rsc_rls_obj_ld_core_sct = dout_8_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_dp
    (
  clk, rst, dout_9_rsc_req_obj_oswt, dout_9_rsc_req_obj_wen_comp, dout_9_rsc_req_obj_biwt,
      dout_9_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_9_rsc_req_obj_oswt;
  output dout_9_rsc_req_obj_wen_comp;
  input dout_9_rsc_req_obj_biwt;
  input dout_9_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_9_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_9_rsc_req_obj_wen_comp = (~ dout_9_rsc_req_obj_oswt) | dout_9_rsc_req_obj_biwt
      | dout_9_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_9_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_9_rsc_req_obj_bcwt <= ~((~(dout_9_rsc_req_obj_bcwt | dout_9_rsc_req_obj_biwt))
          | dout_9_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_9_rsc_req_obj_oswt, dout_9_rsc_req_obj_vd,
      dout_9_rsc_req_obj_biwt, dout_9_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_9_rsc_req_obj_oswt;
  input dout_9_rsc_req_obj_vd;
  output dout_9_rsc_req_obj_biwt;
  output dout_9_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_9_rsc_req_obj_pdswt0;
  reg dout_9_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_9_rsc_req_obj_pdswt0 = (~ core_wten) & dout_9_rsc_req_obj_oswt;
  assign dout_9_rsc_req_obj_biwt = (dout_9_rsc_req_obj_pdswt0 | dout_9_rsc_req_obj_icwt)
      & dout_9_rsc_req_obj_vd;
  assign dout_9_rsc_req_obj_bdwt = dout_9_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_9_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_9_rsc_req_obj_icwt <= ~((~(dout_9_rsc_req_obj_icwt | dout_9_rsc_req_obj_pdswt0))
          | dout_9_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_rls_obj_dout_9_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_rls_obj_dout_9_rsc_rls_wait_ctrl
    (
  core_wten, dout_9_rsc_rls_obj_iswt0, dout_9_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_9_rsc_rls_obj_iswt0;
  output dout_9_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_9_rsc_rls_obj_ld_core_sct = dout_9_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_dp
    (
  clk, rst, dout_10_rsc_req_obj_oswt, dout_10_rsc_req_obj_wen_comp, dout_10_rsc_req_obj_biwt,
      dout_10_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_10_rsc_req_obj_oswt;
  output dout_10_rsc_req_obj_wen_comp;
  input dout_10_rsc_req_obj_biwt;
  input dout_10_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_10_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_10_rsc_req_obj_wen_comp = (~ dout_10_rsc_req_obj_oswt) | dout_10_rsc_req_obj_biwt
      | dout_10_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_10_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_10_rsc_req_obj_bcwt <= ~((~(dout_10_rsc_req_obj_bcwt | dout_10_rsc_req_obj_biwt))
          | dout_10_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_10_rsc_req_obj_oswt, dout_10_rsc_req_obj_vd,
      dout_10_rsc_req_obj_biwt, dout_10_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_10_rsc_req_obj_oswt;
  input dout_10_rsc_req_obj_vd;
  output dout_10_rsc_req_obj_biwt;
  output dout_10_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_10_rsc_req_obj_pdswt0;
  reg dout_10_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_10_rsc_req_obj_pdswt0 = (~ core_wten) & dout_10_rsc_req_obj_oswt;
  assign dout_10_rsc_req_obj_biwt = (dout_10_rsc_req_obj_pdswt0 | dout_10_rsc_req_obj_icwt)
      & dout_10_rsc_req_obj_vd;
  assign dout_10_rsc_req_obj_bdwt = dout_10_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_10_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_10_rsc_req_obj_icwt <= ~((~(dout_10_rsc_req_obj_icwt | dout_10_rsc_req_obj_pdswt0))
          | dout_10_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_rls_obj_dout_10_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_rls_obj_dout_10_rsc_rls_wait_ctrl
    (
  core_wten, dout_10_rsc_rls_obj_iswt0, dout_10_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_10_rsc_rls_obj_iswt0;
  output dout_10_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_10_rsc_rls_obj_ld_core_sct = dout_10_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_dp
    (
  clk, rst, dout_11_rsc_req_obj_oswt, dout_11_rsc_req_obj_wen_comp, dout_11_rsc_req_obj_biwt,
      dout_11_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_11_rsc_req_obj_oswt;
  output dout_11_rsc_req_obj_wen_comp;
  input dout_11_rsc_req_obj_biwt;
  input dout_11_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_11_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_11_rsc_req_obj_wen_comp = (~ dout_11_rsc_req_obj_oswt) | dout_11_rsc_req_obj_biwt
      | dout_11_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_11_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_11_rsc_req_obj_bcwt <= ~((~(dout_11_rsc_req_obj_bcwt | dout_11_rsc_req_obj_biwt))
          | dout_11_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_11_rsc_req_obj_oswt, dout_11_rsc_req_obj_vd,
      dout_11_rsc_req_obj_biwt, dout_11_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_11_rsc_req_obj_oswt;
  input dout_11_rsc_req_obj_vd;
  output dout_11_rsc_req_obj_biwt;
  output dout_11_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_11_rsc_req_obj_pdswt0;
  reg dout_11_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_11_rsc_req_obj_pdswt0 = (~ core_wten) & dout_11_rsc_req_obj_oswt;
  assign dout_11_rsc_req_obj_biwt = (dout_11_rsc_req_obj_pdswt0 | dout_11_rsc_req_obj_icwt)
      & dout_11_rsc_req_obj_vd;
  assign dout_11_rsc_req_obj_bdwt = dout_11_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_11_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_11_rsc_req_obj_icwt <= ~((~(dout_11_rsc_req_obj_icwt | dout_11_rsc_req_obj_pdswt0))
          | dout_11_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_rls_obj_dout_11_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_rls_obj_dout_11_rsc_rls_wait_ctrl
    (
  core_wten, dout_11_rsc_rls_obj_iswt0, dout_11_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_11_rsc_rls_obj_iswt0;
  output dout_11_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_11_rsc_rls_obj_ld_core_sct = dout_11_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_dp
    (
  clk, rst, dout_12_rsc_req_obj_oswt, dout_12_rsc_req_obj_wen_comp, dout_12_rsc_req_obj_biwt,
      dout_12_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_12_rsc_req_obj_oswt;
  output dout_12_rsc_req_obj_wen_comp;
  input dout_12_rsc_req_obj_biwt;
  input dout_12_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_12_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_12_rsc_req_obj_wen_comp = (~ dout_12_rsc_req_obj_oswt) | dout_12_rsc_req_obj_biwt
      | dout_12_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_12_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_12_rsc_req_obj_bcwt <= ~((~(dout_12_rsc_req_obj_bcwt | dout_12_rsc_req_obj_biwt))
          | dout_12_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_12_rsc_req_obj_oswt, dout_12_rsc_req_obj_vd,
      dout_12_rsc_req_obj_biwt, dout_12_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_12_rsc_req_obj_oswt;
  input dout_12_rsc_req_obj_vd;
  output dout_12_rsc_req_obj_biwt;
  output dout_12_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_12_rsc_req_obj_pdswt0;
  reg dout_12_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_12_rsc_req_obj_pdswt0 = (~ core_wten) & dout_12_rsc_req_obj_oswt;
  assign dout_12_rsc_req_obj_biwt = (dout_12_rsc_req_obj_pdswt0 | dout_12_rsc_req_obj_icwt)
      & dout_12_rsc_req_obj_vd;
  assign dout_12_rsc_req_obj_bdwt = dout_12_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_12_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_12_rsc_req_obj_icwt <= ~((~(dout_12_rsc_req_obj_icwt | dout_12_rsc_req_obj_pdswt0))
          | dout_12_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_rls_obj_dout_12_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_rls_obj_dout_12_rsc_rls_wait_ctrl
    (
  core_wten, dout_12_rsc_rls_obj_iswt0, dout_12_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_12_rsc_rls_obj_iswt0;
  output dout_12_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_12_rsc_rls_obj_ld_core_sct = dout_12_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_dp
    (
  clk, rst, dout_13_rsc_req_obj_oswt, dout_13_rsc_req_obj_wen_comp, dout_13_rsc_req_obj_biwt,
      dout_13_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_13_rsc_req_obj_oswt;
  output dout_13_rsc_req_obj_wen_comp;
  input dout_13_rsc_req_obj_biwt;
  input dout_13_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_13_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_13_rsc_req_obj_wen_comp = (~ dout_13_rsc_req_obj_oswt) | dout_13_rsc_req_obj_biwt
      | dout_13_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_13_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_13_rsc_req_obj_bcwt <= ~((~(dout_13_rsc_req_obj_bcwt | dout_13_rsc_req_obj_biwt))
          | dout_13_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_13_rsc_req_obj_oswt, dout_13_rsc_req_obj_vd,
      dout_13_rsc_req_obj_biwt, dout_13_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_13_rsc_req_obj_oswt;
  input dout_13_rsc_req_obj_vd;
  output dout_13_rsc_req_obj_biwt;
  output dout_13_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_13_rsc_req_obj_pdswt0;
  reg dout_13_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_13_rsc_req_obj_pdswt0 = (~ core_wten) & dout_13_rsc_req_obj_oswt;
  assign dout_13_rsc_req_obj_biwt = (dout_13_rsc_req_obj_pdswt0 | dout_13_rsc_req_obj_icwt)
      & dout_13_rsc_req_obj_vd;
  assign dout_13_rsc_req_obj_bdwt = dout_13_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_13_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_13_rsc_req_obj_icwt <= ~((~(dout_13_rsc_req_obj_icwt | dout_13_rsc_req_obj_pdswt0))
          | dout_13_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_rls_obj_dout_13_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_rls_obj_dout_13_rsc_rls_wait_ctrl
    (
  core_wten, dout_13_rsc_rls_obj_iswt0, dout_13_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_13_rsc_rls_obj_iswt0;
  output dout_13_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_13_rsc_rls_obj_ld_core_sct = dout_13_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_dp
    (
  clk, rst, dout_14_rsc_req_obj_oswt, dout_14_rsc_req_obj_wen_comp, dout_14_rsc_req_obj_biwt,
      dout_14_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_14_rsc_req_obj_oswt;
  output dout_14_rsc_req_obj_wen_comp;
  input dout_14_rsc_req_obj_biwt;
  input dout_14_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_14_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_14_rsc_req_obj_wen_comp = (~ dout_14_rsc_req_obj_oswt) | dout_14_rsc_req_obj_biwt
      | dout_14_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_14_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_14_rsc_req_obj_bcwt <= ~((~(dout_14_rsc_req_obj_bcwt | dout_14_rsc_req_obj_biwt))
          | dout_14_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_14_rsc_req_obj_oswt, dout_14_rsc_req_obj_vd,
      dout_14_rsc_req_obj_biwt, dout_14_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_14_rsc_req_obj_oswt;
  input dout_14_rsc_req_obj_vd;
  output dout_14_rsc_req_obj_biwt;
  output dout_14_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_14_rsc_req_obj_pdswt0;
  reg dout_14_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_14_rsc_req_obj_pdswt0 = (~ core_wten) & dout_14_rsc_req_obj_oswt;
  assign dout_14_rsc_req_obj_biwt = (dout_14_rsc_req_obj_pdswt0 | dout_14_rsc_req_obj_icwt)
      & dout_14_rsc_req_obj_vd;
  assign dout_14_rsc_req_obj_bdwt = dout_14_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_14_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_14_rsc_req_obj_icwt <= ~((~(dout_14_rsc_req_obj_icwt | dout_14_rsc_req_obj_pdswt0))
          | dout_14_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_rls_obj_dout_14_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_rls_obj_dout_14_rsc_rls_wait_ctrl
    (
  core_wten, dout_14_rsc_rls_obj_iswt0, dout_14_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_14_rsc_rls_obj_iswt0;
  output dout_14_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_14_rsc_rls_obj_ld_core_sct = dout_14_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_dp
    (
  clk, rst, dout_15_rsc_req_obj_oswt, dout_15_rsc_req_obj_wen_comp, dout_15_rsc_req_obj_biwt,
      dout_15_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_15_rsc_req_obj_oswt;
  output dout_15_rsc_req_obj_wen_comp;
  input dout_15_rsc_req_obj_biwt;
  input dout_15_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_15_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_15_rsc_req_obj_wen_comp = (~ dout_15_rsc_req_obj_oswt) | dout_15_rsc_req_obj_biwt
      | dout_15_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_15_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_15_rsc_req_obj_bcwt <= ~((~(dout_15_rsc_req_obj_bcwt | dout_15_rsc_req_obj_biwt))
          | dout_15_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_15_rsc_req_obj_oswt, dout_15_rsc_req_obj_vd,
      dout_15_rsc_req_obj_biwt, dout_15_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_15_rsc_req_obj_oswt;
  input dout_15_rsc_req_obj_vd;
  output dout_15_rsc_req_obj_biwt;
  output dout_15_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_15_rsc_req_obj_pdswt0;
  reg dout_15_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_15_rsc_req_obj_pdswt0 = (~ core_wten) & dout_15_rsc_req_obj_oswt;
  assign dout_15_rsc_req_obj_biwt = (dout_15_rsc_req_obj_pdswt0 | dout_15_rsc_req_obj_icwt)
      & dout_15_rsc_req_obj_vd;
  assign dout_15_rsc_req_obj_bdwt = dout_15_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_15_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_15_rsc_req_obj_icwt <= ~((~(dout_15_rsc_req_obj_icwt | dout_15_rsc_req_obj_pdswt0))
          | dout_15_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_rls_obj_dout_15_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_rls_obj_dout_15_rsc_rls_wait_ctrl
    (
  core_wten, dout_15_rsc_rls_obj_iswt0, dout_15_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_15_rsc_rls_obj_iswt0;
  output dout_15_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_15_rsc_rls_obj_ld_core_sct = dout_15_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj_dout_16_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj_dout_16_rsc_req_wait_dp
    (
  clk, rst, dout_16_rsc_req_obj_oswt, dout_16_rsc_req_obj_wen_comp, dout_16_rsc_req_obj_biwt,
      dout_16_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_16_rsc_req_obj_oswt;
  output dout_16_rsc_req_obj_wen_comp;
  input dout_16_rsc_req_obj_biwt;
  input dout_16_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_16_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_16_rsc_req_obj_wen_comp = (~ dout_16_rsc_req_obj_oswt) | dout_16_rsc_req_obj_biwt
      | dout_16_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_16_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_16_rsc_req_obj_bcwt <= ~((~(dout_16_rsc_req_obj_bcwt | dout_16_rsc_req_obj_biwt))
          | dout_16_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj_dout_16_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj_dout_16_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_16_rsc_req_obj_oswt, dout_16_rsc_req_obj_vd,
      dout_16_rsc_req_obj_biwt, dout_16_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_16_rsc_req_obj_oswt;
  input dout_16_rsc_req_obj_vd;
  output dout_16_rsc_req_obj_biwt;
  output dout_16_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_16_rsc_req_obj_pdswt0;
  reg dout_16_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_16_rsc_req_obj_pdswt0 = (~ core_wten) & dout_16_rsc_req_obj_oswt;
  assign dout_16_rsc_req_obj_biwt = (dout_16_rsc_req_obj_pdswt0 | dout_16_rsc_req_obj_icwt)
      & dout_16_rsc_req_obj_vd;
  assign dout_16_rsc_req_obj_bdwt = dout_16_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_16_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_16_rsc_req_obj_icwt <= ~((~(dout_16_rsc_req_obj_icwt | dout_16_rsc_req_obj_pdswt0))
          | dout_16_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_rls_obj_dout_16_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_rls_obj_dout_16_rsc_rls_wait_ctrl
    (
  core_wten, dout_16_rsc_rls_obj_iswt0, dout_16_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_16_rsc_rls_obj_iswt0;
  output dout_16_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_16_rsc_rls_obj_ld_core_sct = dout_16_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj_dout_17_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj_dout_17_rsc_req_wait_dp
    (
  clk, rst, dout_17_rsc_req_obj_oswt, dout_17_rsc_req_obj_wen_comp, dout_17_rsc_req_obj_biwt,
      dout_17_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_17_rsc_req_obj_oswt;
  output dout_17_rsc_req_obj_wen_comp;
  input dout_17_rsc_req_obj_biwt;
  input dout_17_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_17_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_17_rsc_req_obj_wen_comp = (~ dout_17_rsc_req_obj_oswt) | dout_17_rsc_req_obj_biwt
      | dout_17_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_17_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_17_rsc_req_obj_bcwt <= ~((~(dout_17_rsc_req_obj_bcwt | dout_17_rsc_req_obj_biwt))
          | dout_17_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj_dout_17_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj_dout_17_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_17_rsc_req_obj_oswt, dout_17_rsc_req_obj_vd,
      dout_17_rsc_req_obj_biwt, dout_17_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_17_rsc_req_obj_oswt;
  input dout_17_rsc_req_obj_vd;
  output dout_17_rsc_req_obj_biwt;
  output dout_17_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_17_rsc_req_obj_pdswt0;
  reg dout_17_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_17_rsc_req_obj_pdswt0 = (~ core_wten) & dout_17_rsc_req_obj_oswt;
  assign dout_17_rsc_req_obj_biwt = (dout_17_rsc_req_obj_pdswt0 | dout_17_rsc_req_obj_icwt)
      & dout_17_rsc_req_obj_vd;
  assign dout_17_rsc_req_obj_bdwt = dout_17_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_17_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_17_rsc_req_obj_icwt <= ~((~(dout_17_rsc_req_obj_icwt | dout_17_rsc_req_obj_pdswt0))
          | dout_17_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_rls_obj_dout_17_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_rls_obj_dout_17_rsc_rls_wait_ctrl
    (
  core_wten, dout_17_rsc_rls_obj_iswt0, dout_17_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_17_rsc_rls_obj_iswt0;
  output dout_17_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_17_rsc_rls_obj_ld_core_sct = dout_17_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_dp
    (
  clk, rst, tmp_17_data_rsci_addra_d, tmp_17_data_rsci_addrb_d, tmp_17_data_rsci_douta_d,
      tmp_17_data_rsci_addra_d_core, tmp_17_data_rsci_addrb_d_core, tmp_17_data_rsci_douta_d_mxwt,
      tmp_17_data_rsci_biwt, tmp_17_data_rsci_bdwt, tmp_17_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_17_data_rsci_addra_d;
  output [7:0] tmp_17_data_rsci_addrb_d;
  input [63:0] tmp_17_data_rsci_douta_d;
  input [7:0] tmp_17_data_rsci_addra_d_core;
  input [7:0] tmp_17_data_rsci_addrb_d_core;
  output [15:0] tmp_17_data_rsci_douta_d_mxwt;
  input tmp_17_data_rsci_biwt;
  input tmp_17_data_rsci_bdwt;
  input tmp_17_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_17_data_rsci_bcwt;
  reg [15:0] tmp_17_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_17_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_17_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_17_data_rsci_douta_d[15:0]),
      tmp_17_data_rsci_douta_d_bfwt_15_0, tmp_17_data_rsci_bcwt);
  assign tmp_17_data_rsci_douta_d_mxwt = tmp_17_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_17_data_rsci_addra_d = {(~ tmp_17_data_rsci_biwt_pff) , (tmp_17_data_rsci_addra_d_core[6:0])};
  assign tmp_17_data_rsci_addrb_d = {(~ tmp_17_data_rsci_biwt_pff) , (tmp_17_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_17_data_rsci_bcwt <= 1'b0;
      tmp_17_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_17_data_rsci_bcwt <= ~((~(tmp_17_data_rsci_bcwt | tmp_17_data_rsci_biwt))
          | tmp_17_data_rsci_bdwt);
      tmp_17_data_rsci_douta_d_bfwt_15_0 <= tmp_17_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_17_data_rsci_oswt, tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_17_data_rsci_biwt,
      tmp_17_data_rsci_bdwt, tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_17_data_rsci_biwt_pff,
      tmp_17_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_17_data_rsci_oswt;
  input tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_17_data_rsci_biwt;
  output tmp_17_data_rsci_bdwt;
  output tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_17_data_rsci_biwt_pff;
  input tmp_17_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_17_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_17_data_rsci_bdwt = tmp_17_data_rsci_oswt & core_wen;
  assign tmp_17_data_rsci_biwt = (~ core_wten) & tmp_17_data_rsci_oswt;
  assign tmp_17_data_rsci_biwt_pff = tmp_17_data_rsci_tiswt0_pff;
  assign tmp_17_data_rsci_tiswt0_pff = core_wen & tmp_17_data_rsci_oswt_pff;
  assign tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_17_data_rsci_tiswt0_pff;
  assign tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_17_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_dp
    (
  clk, rst, tmp_16_data_rsci_addra_d, tmp_16_data_rsci_addrb_d, tmp_16_data_rsci_douta_d,
      tmp_16_data_rsci_addra_d_core, tmp_16_data_rsci_addrb_d_core, tmp_16_data_rsci_douta_d_mxwt,
      tmp_16_data_rsci_biwt, tmp_16_data_rsci_bdwt, tmp_16_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_16_data_rsci_addra_d;
  output [7:0] tmp_16_data_rsci_addrb_d;
  input [63:0] tmp_16_data_rsci_douta_d;
  input [7:0] tmp_16_data_rsci_addra_d_core;
  input [7:0] tmp_16_data_rsci_addrb_d_core;
  output [15:0] tmp_16_data_rsci_douta_d_mxwt;
  input tmp_16_data_rsci_biwt;
  input tmp_16_data_rsci_bdwt;
  input tmp_16_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_16_data_rsci_bcwt;
  reg [15:0] tmp_16_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_16_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_16_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_16_data_rsci_douta_d[15:0]),
      tmp_16_data_rsci_douta_d_bfwt_15_0, tmp_16_data_rsci_bcwt);
  assign tmp_16_data_rsci_douta_d_mxwt = tmp_16_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_16_data_rsci_addra_d = {(~ tmp_16_data_rsci_biwt_pff) , (tmp_16_data_rsci_addra_d_core[6:0])};
  assign tmp_16_data_rsci_addrb_d = {(~ tmp_16_data_rsci_biwt_pff) , (tmp_16_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_16_data_rsci_bcwt <= 1'b0;
      tmp_16_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_16_data_rsci_bcwt <= ~((~(tmp_16_data_rsci_bcwt | tmp_16_data_rsci_biwt))
          | tmp_16_data_rsci_bdwt);
      tmp_16_data_rsci_douta_d_bfwt_15_0 <= tmp_16_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_16_data_rsci_oswt, tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_16_data_rsci_biwt,
      tmp_16_data_rsci_bdwt, tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_16_data_rsci_biwt_pff,
      tmp_16_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_16_data_rsci_oswt;
  input tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_16_data_rsci_biwt;
  output tmp_16_data_rsci_bdwt;
  output tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_16_data_rsci_biwt_pff;
  input tmp_16_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_16_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_16_data_rsci_bdwt = tmp_16_data_rsci_oswt & core_wen;
  assign tmp_16_data_rsci_biwt = (~ core_wten) & tmp_16_data_rsci_oswt;
  assign tmp_16_data_rsci_biwt_pff = tmp_16_data_rsci_tiswt0_pff;
  assign tmp_16_data_rsci_tiswt0_pff = core_wen & tmp_16_data_rsci_oswt_pff;
  assign tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_16_data_rsci_tiswt0_pff;
  assign tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_16_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_dp
    (
  clk, rst, tmp_15_data_rsci_addra_d, tmp_15_data_rsci_addrb_d, tmp_15_data_rsci_douta_d,
      tmp_15_data_rsci_addra_d_core, tmp_15_data_rsci_addrb_d_core, tmp_15_data_rsci_douta_d_mxwt,
      tmp_15_data_rsci_biwt, tmp_15_data_rsci_bdwt, tmp_15_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_15_data_rsci_addra_d;
  output [7:0] tmp_15_data_rsci_addrb_d;
  input [63:0] tmp_15_data_rsci_douta_d;
  input [7:0] tmp_15_data_rsci_addra_d_core;
  input [7:0] tmp_15_data_rsci_addrb_d_core;
  output [15:0] tmp_15_data_rsci_douta_d_mxwt;
  input tmp_15_data_rsci_biwt;
  input tmp_15_data_rsci_bdwt;
  input tmp_15_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_15_data_rsci_bcwt;
  reg [15:0] tmp_15_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_15_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_15_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_15_data_rsci_douta_d[15:0]),
      tmp_15_data_rsci_douta_d_bfwt_15_0, tmp_15_data_rsci_bcwt);
  assign tmp_15_data_rsci_douta_d_mxwt = tmp_15_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_15_data_rsci_addra_d = {(~ tmp_15_data_rsci_biwt_pff) , (tmp_15_data_rsci_addra_d_core[6:0])};
  assign tmp_15_data_rsci_addrb_d = {(~ tmp_15_data_rsci_biwt_pff) , (tmp_15_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_15_data_rsci_bcwt <= 1'b0;
      tmp_15_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_15_data_rsci_bcwt <= ~((~(tmp_15_data_rsci_bcwt | tmp_15_data_rsci_biwt))
          | tmp_15_data_rsci_bdwt);
      tmp_15_data_rsci_douta_d_bfwt_15_0 <= tmp_15_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_15_data_rsci_oswt, tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_15_data_rsci_biwt,
      tmp_15_data_rsci_bdwt, tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_15_data_rsci_biwt_pff,
      tmp_15_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_15_data_rsci_oswt;
  input tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_15_data_rsci_biwt;
  output tmp_15_data_rsci_bdwt;
  output tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_15_data_rsci_biwt_pff;
  input tmp_15_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_15_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_15_data_rsci_bdwt = tmp_15_data_rsci_oswt & core_wen;
  assign tmp_15_data_rsci_biwt = (~ core_wten) & tmp_15_data_rsci_oswt;
  assign tmp_15_data_rsci_biwt_pff = tmp_15_data_rsci_tiswt0_pff;
  assign tmp_15_data_rsci_tiswt0_pff = core_wen & tmp_15_data_rsci_oswt_pff;
  assign tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_15_data_rsci_tiswt0_pff;
  assign tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_15_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_dp
    (
  clk, rst, tmp_14_data_rsci_addra_d, tmp_14_data_rsci_addrb_d, tmp_14_data_rsci_douta_d,
      tmp_14_data_rsci_addra_d_core, tmp_14_data_rsci_addrb_d_core, tmp_14_data_rsci_douta_d_mxwt,
      tmp_14_data_rsci_biwt, tmp_14_data_rsci_bdwt, tmp_14_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_14_data_rsci_addra_d;
  output [7:0] tmp_14_data_rsci_addrb_d;
  input [63:0] tmp_14_data_rsci_douta_d;
  input [7:0] tmp_14_data_rsci_addra_d_core;
  input [7:0] tmp_14_data_rsci_addrb_d_core;
  output [15:0] tmp_14_data_rsci_douta_d_mxwt;
  input tmp_14_data_rsci_biwt;
  input tmp_14_data_rsci_bdwt;
  input tmp_14_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_14_data_rsci_bcwt;
  reg [15:0] tmp_14_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_14_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_14_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_14_data_rsci_douta_d[15:0]),
      tmp_14_data_rsci_douta_d_bfwt_15_0, tmp_14_data_rsci_bcwt);
  assign tmp_14_data_rsci_douta_d_mxwt = tmp_14_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_14_data_rsci_addra_d = {(~ tmp_14_data_rsci_biwt_pff) , (tmp_14_data_rsci_addra_d_core[6:0])};
  assign tmp_14_data_rsci_addrb_d = {(~ tmp_14_data_rsci_biwt_pff) , (tmp_14_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_14_data_rsci_bcwt <= 1'b0;
      tmp_14_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_14_data_rsci_bcwt <= ~((~(tmp_14_data_rsci_bcwt | tmp_14_data_rsci_biwt))
          | tmp_14_data_rsci_bdwt);
      tmp_14_data_rsci_douta_d_bfwt_15_0 <= tmp_14_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_14_data_rsci_oswt, tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_14_data_rsci_biwt,
      tmp_14_data_rsci_bdwt, tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_14_data_rsci_biwt_pff,
      tmp_14_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_14_data_rsci_oswt;
  input tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_14_data_rsci_biwt;
  output tmp_14_data_rsci_bdwt;
  output tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_14_data_rsci_biwt_pff;
  input tmp_14_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_14_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_14_data_rsci_bdwt = tmp_14_data_rsci_oswt & core_wen;
  assign tmp_14_data_rsci_biwt = (~ core_wten) & tmp_14_data_rsci_oswt;
  assign tmp_14_data_rsci_biwt_pff = tmp_14_data_rsci_tiswt0_pff;
  assign tmp_14_data_rsci_tiswt0_pff = core_wen & tmp_14_data_rsci_oswt_pff;
  assign tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_14_data_rsci_tiswt0_pff;
  assign tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_14_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_dp
    (
  clk, rst, tmp_13_data_rsci_addra_d, tmp_13_data_rsci_addrb_d, tmp_13_data_rsci_douta_d,
      tmp_13_data_rsci_addra_d_core, tmp_13_data_rsci_addrb_d_core, tmp_13_data_rsci_douta_d_mxwt,
      tmp_13_data_rsci_biwt, tmp_13_data_rsci_bdwt, tmp_13_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_13_data_rsci_addra_d;
  output [7:0] tmp_13_data_rsci_addrb_d;
  input [63:0] tmp_13_data_rsci_douta_d;
  input [7:0] tmp_13_data_rsci_addra_d_core;
  input [7:0] tmp_13_data_rsci_addrb_d_core;
  output [15:0] tmp_13_data_rsci_douta_d_mxwt;
  input tmp_13_data_rsci_biwt;
  input tmp_13_data_rsci_bdwt;
  input tmp_13_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_13_data_rsci_bcwt;
  reg [15:0] tmp_13_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_13_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_13_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_13_data_rsci_douta_d[15:0]),
      tmp_13_data_rsci_douta_d_bfwt_15_0, tmp_13_data_rsci_bcwt);
  assign tmp_13_data_rsci_douta_d_mxwt = tmp_13_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_13_data_rsci_addra_d = {(~ tmp_13_data_rsci_biwt_pff) , (tmp_13_data_rsci_addra_d_core[6:0])};
  assign tmp_13_data_rsci_addrb_d = {(~ tmp_13_data_rsci_biwt_pff) , (tmp_13_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_13_data_rsci_bcwt <= 1'b0;
      tmp_13_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_13_data_rsci_bcwt <= ~((~(tmp_13_data_rsci_bcwt | tmp_13_data_rsci_biwt))
          | tmp_13_data_rsci_bdwt);
      tmp_13_data_rsci_douta_d_bfwt_15_0 <= tmp_13_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_13_data_rsci_oswt, tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_13_data_rsci_biwt,
      tmp_13_data_rsci_bdwt, tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_13_data_rsci_biwt_pff,
      tmp_13_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_13_data_rsci_oswt;
  input tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_13_data_rsci_biwt;
  output tmp_13_data_rsci_bdwt;
  output tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_13_data_rsci_biwt_pff;
  input tmp_13_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_13_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_13_data_rsci_bdwt = tmp_13_data_rsci_oswt & core_wen;
  assign tmp_13_data_rsci_biwt = (~ core_wten) & tmp_13_data_rsci_oswt;
  assign tmp_13_data_rsci_biwt_pff = tmp_13_data_rsci_tiswt0_pff;
  assign tmp_13_data_rsci_tiswt0_pff = core_wen & tmp_13_data_rsci_oswt_pff;
  assign tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_13_data_rsci_tiswt0_pff;
  assign tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_13_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_dp
    (
  clk, rst, tmp_12_data_rsci_addra_d, tmp_12_data_rsci_addrb_d, tmp_12_data_rsci_douta_d,
      tmp_12_data_rsci_addra_d_core, tmp_12_data_rsci_addrb_d_core, tmp_12_data_rsci_douta_d_mxwt,
      tmp_12_data_rsci_biwt, tmp_12_data_rsci_bdwt, tmp_12_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_12_data_rsci_addra_d;
  output [7:0] tmp_12_data_rsci_addrb_d;
  input [63:0] tmp_12_data_rsci_douta_d;
  input [7:0] tmp_12_data_rsci_addra_d_core;
  input [7:0] tmp_12_data_rsci_addrb_d_core;
  output [15:0] tmp_12_data_rsci_douta_d_mxwt;
  input tmp_12_data_rsci_biwt;
  input tmp_12_data_rsci_bdwt;
  input tmp_12_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_12_data_rsci_bcwt;
  reg [15:0] tmp_12_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_12_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_12_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_12_data_rsci_douta_d[15:0]),
      tmp_12_data_rsci_douta_d_bfwt_15_0, tmp_12_data_rsci_bcwt);
  assign tmp_12_data_rsci_douta_d_mxwt = tmp_12_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_12_data_rsci_addra_d = {(~ tmp_12_data_rsci_biwt_pff) , (tmp_12_data_rsci_addra_d_core[6:0])};
  assign tmp_12_data_rsci_addrb_d = {(~ tmp_12_data_rsci_biwt_pff) , (tmp_12_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_12_data_rsci_bcwt <= 1'b0;
      tmp_12_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_12_data_rsci_bcwt <= ~((~(tmp_12_data_rsci_bcwt | tmp_12_data_rsci_biwt))
          | tmp_12_data_rsci_bdwt);
      tmp_12_data_rsci_douta_d_bfwt_15_0 <= tmp_12_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_12_data_rsci_oswt, tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_12_data_rsci_biwt,
      tmp_12_data_rsci_bdwt, tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_12_data_rsci_biwt_pff,
      tmp_12_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_12_data_rsci_oswt;
  input tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_12_data_rsci_biwt;
  output tmp_12_data_rsci_bdwt;
  output tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_12_data_rsci_biwt_pff;
  input tmp_12_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_12_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_12_data_rsci_bdwt = tmp_12_data_rsci_oswt & core_wen;
  assign tmp_12_data_rsci_biwt = (~ core_wten) & tmp_12_data_rsci_oswt;
  assign tmp_12_data_rsci_biwt_pff = tmp_12_data_rsci_tiswt0_pff;
  assign tmp_12_data_rsci_tiswt0_pff = core_wen & tmp_12_data_rsci_oswt_pff;
  assign tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_12_data_rsci_tiswt0_pff;
  assign tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_12_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_dp
    (
  clk, rst, tmp_11_data_rsci_addra_d, tmp_11_data_rsci_addrb_d, tmp_11_data_rsci_douta_d,
      tmp_11_data_rsci_addra_d_core, tmp_11_data_rsci_addrb_d_core, tmp_11_data_rsci_douta_d_mxwt,
      tmp_11_data_rsci_biwt, tmp_11_data_rsci_bdwt, tmp_11_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_11_data_rsci_addra_d;
  output [7:0] tmp_11_data_rsci_addrb_d;
  input [63:0] tmp_11_data_rsci_douta_d;
  input [7:0] tmp_11_data_rsci_addra_d_core;
  input [7:0] tmp_11_data_rsci_addrb_d_core;
  output [15:0] tmp_11_data_rsci_douta_d_mxwt;
  input tmp_11_data_rsci_biwt;
  input tmp_11_data_rsci_bdwt;
  input tmp_11_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_11_data_rsci_bcwt;
  reg [15:0] tmp_11_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_11_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_11_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_11_data_rsci_douta_d[15:0]),
      tmp_11_data_rsci_douta_d_bfwt_15_0, tmp_11_data_rsci_bcwt);
  assign tmp_11_data_rsci_douta_d_mxwt = tmp_11_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_11_data_rsci_addra_d = {(~ tmp_11_data_rsci_biwt_pff) , (tmp_11_data_rsci_addra_d_core[6:0])};
  assign tmp_11_data_rsci_addrb_d = {(~ tmp_11_data_rsci_biwt_pff) , (tmp_11_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_11_data_rsci_bcwt <= 1'b0;
      tmp_11_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_11_data_rsci_bcwt <= ~((~(tmp_11_data_rsci_bcwt | tmp_11_data_rsci_biwt))
          | tmp_11_data_rsci_bdwt);
      tmp_11_data_rsci_douta_d_bfwt_15_0 <= tmp_11_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_11_data_rsci_oswt, tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_11_data_rsci_biwt,
      tmp_11_data_rsci_bdwt, tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_11_data_rsci_biwt_pff,
      tmp_11_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_11_data_rsci_oswt;
  input tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_11_data_rsci_biwt;
  output tmp_11_data_rsci_bdwt;
  output tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_11_data_rsci_biwt_pff;
  input tmp_11_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_11_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_11_data_rsci_bdwt = tmp_11_data_rsci_oswt & core_wen;
  assign tmp_11_data_rsci_biwt = (~ core_wten) & tmp_11_data_rsci_oswt;
  assign tmp_11_data_rsci_biwt_pff = tmp_11_data_rsci_tiswt0_pff;
  assign tmp_11_data_rsci_tiswt0_pff = core_wen & tmp_11_data_rsci_oswt_pff;
  assign tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_11_data_rsci_tiswt0_pff;
  assign tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_11_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_dp
    (
  clk, rst, tmp_10_data_rsci_addra_d, tmp_10_data_rsci_addrb_d, tmp_10_data_rsci_douta_d,
      tmp_10_data_rsci_addra_d_core, tmp_10_data_rsci_addrb_d_core, tmp_10_data_rsci_douta_d_mxwt,
      tmp_10_data_rsci_biwt, tmp_10_data_rsci_bdwt, tmp_10_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_10_data_rsci_addra_d;
  output [7:0] tmp_10_data_rsci_addrb_d;
  input [63:0] tmp_10_data_rsci_douta_d;
  input [7:0] tmp_10_data_rsci_addra_d_core;
  input [7:0] tmp_10_data_rsci_addrb_d_core;
  output [15:0] tmp_10_data_rsci_douta_d_mxwt;
  input tmp_10_data_rsci_biwt;
  input tmp_10_data_rsci_bdwt;
  input tmp_10_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_10_data_rsci_bcwt;
  reg [15:0] tmp_10_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_10_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_10_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_10_data_rsci_douta_d[15:0]),
      tmp_10_data_rsci_douta_d_bfwt_15_0, tmp_10_data_rsci_bcwt);
  assign tmp_10_data_rsci_douta_d_mxwt = tmp_10_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_10_data_rsci_addra_d = {(~ tmp_10_data_rsci_biwt_pff) , (tmp_10_data_rsci_addra_d_core[6:0])};
  assign tmp_10_data_rsci_addrb_d = {(~ tmp_10_data_rsci_biwt_pff) , (tmp_10_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_10_data_rsci_bcwt <= 1'b0;
      tmp_10_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_10_data_rsci_bcwt <= ~((~(tmp_10_data_rsci_bcwt | tmp_10_data_rsci_biwt))
          | tmp_10_data_rsci_bdwt);
      tmp_10_data_rsci_douta_d_bfwt_15_0 <= tmp_10_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_10_data_rsci_oswt, tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_10_data_rsci_biwt,
      tmp_10_data_rsci_bdwt, tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_10_data_rsci_biwt_pff,
      tmp_10_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_10_data_rsci_oswt;
  input tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_10_data_rsci_biwt;
  output tmp_10_data_rsci_bdwt;
  output tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_10_data_rsci_biwt_pff;
  input tmp_10_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_10_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_10_data_rsci_bdwt = tmp_10_data_rsci_oswt & core_wen;
  assign tmp_10_data_rsci_biwt = (~ core_wten) & tmp_10_data_rsci_oswt;
  assign tmp_10_data_rsci_biwt_pff = tmp_10_data_rsci_tiswt0_pff;
  assign tmp_10_data_rsci_tiswt0_pff = core_wen & tmp_10_data_rsci_oswt_pff;
  assign tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_10_data_rsci_tiswt0_pff;
  assign tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_10_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_dp
    (
  clk, rst, tmp_9_data_rsci_addra_d, tmp_9_data_rsci_addrb_d, tmp_9_data_rsci_douta_d,
      tmp_9_data_rsci_addra_d_core, tmp_9_data_rsci_addrb_d_core, tmp_9_data_rsci_douta_d_mxwt,
      tmp_9_data_rsci_biwt, tmp_9_data_rsci_bdwt, tmp_9_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_9_data_rsci_addra_d;
  output [7:0] tmp_9_data_rsci_addrb_d;
  input [63:0] tmp_9_data_rsci_douta_d;
  input [7:0] tmp_9_data_rsci_addra_d_core;
  input [7:0] tmp_9_data_rsci_addrb_d_core;
  output [15:0] tmp_9_data_rsci_douta_d_mxwt;
  input tmp_9_data_rsci_biwt;
  input tmp_9_data_rsci_bdwt;
  input tmp_9_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_9_data_rsci_bcwt;
  reg [15:0] tmp_9_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_9_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_9_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_9_data_rsci_douta_d[15:0]),
      tmp_9_data_rsci_douta_d_bfwt_15_0, tmp_9_data_rsci_bcwt);
  assign tmp_9_data_rsci_douta_d_mxwt = tmp_9_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_9_data_rsci_addra_d = {(~ tmp_9_data_rsci_biwt_pff) , (tmp_9_data_rsci_addra_d_core[6:0])};
  assign tmp_9_data_rsci_addrb_d = {(~ tmp_9_data_rsci_biwt_pff) , (tmp_9_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_9_data_rsci_bcwt <= 1'b0;
      tmp_9_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_9_data_rsci_bcwt <= ~((~(tmp_9_data_rsci_bcwt | tmp_9_data_rsci_biwt))
          | tmp_9_data_rsci_bdwt);
      tmp_9_data_rsci_douta_d_bfwt_15_0 <= tmp_9_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_9_data_rsci_oswt, tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_9_data_rsci_biwt,
      tmp_9_data_rsci_bdwt, tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_9_data_rsci_biwt_pff,
      tmp_9_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_9_data_rsci_oswt;
  input tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_9_data_rsci_biwt;
  output tmp_9_data_rsci_bdwt;
  output tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_9_data_rsci_biwt_pff;
  input tmp_9_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_9_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_9_data_rsci_bdwt = tmp_9_data_rsci_oswt & core_wen;
  assign tmp_9_data_rsci_biwt = (~ core_wten) & tmp_9_data_rsci_oswt;
  assign tmp_9_data_rsci_biwt_pff = tmp_9_data_rsci_tiswt0_pff;
  assign tmp_9_data_rsci_tiswt0_pff = core_wen & tmp_9_data_rsci_oswt_pff;
  assign tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_9_data_rsci_tiswt0_pff;
  assign tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_9_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_dp
    (
  clk, rst, tmp_8_data_rsci_addra_d, tmp_8_data_rsci_addrb_d, tmp_8_data_rsci_douta_d,
      tmp_8_data_rsci_addra_d_core, tmp_8_data_rsci_addrb_d_core, tmp_8_data_rsci_douta_d_mxwt,
      tmp_8_data_rsci_biwt, tmp_8_data_rsci_bdwt, tmp_8_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_8_data_rsci_addra_d;
  output [7:0] tmp_8_data_rsci_addrb_d;
  input [63:0] tmp_8_data_rsci_douta_d;
  input [7:0] tmp_8_data_rsci_addra_d_core;
  input [7:0] tmp_8_data_rsci_addrb_d_core;
  output [15:0] tmp_8_data_rsci_douta_d_mxwt;
  input tmp_8_data_rsci_biwt;
  input tmp_8_data_rsci_bdwt;
  input tmp_8_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_8_data_rsci_bcwt;
  reg [15:0] tmp_8_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_8_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_8_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_8_data_rsci_douta_d[15:0]),
      tmp_8_data_rsci_douta_d_bfwt_15_0, tmp_8_data_rsci_bcwt);
  assign tmp_8_data_rsci_douta_d_mxwt = tmp_8_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_8_data_rsci_addra_d = {(~ tmp_8_data_rsci_biwt_pff) , (tmp_8_data_rsci_addra_d_core[6:0])};
  assign tmp_8_data_rsci_addrb_d = {(~ tmp_8_data_rsci_biwt_pff) , (tmp_8_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_8_data_rsci_bcwt <= 1'b0;
      tmp_8_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_8_data_rsci_bcwt <= ~((~(tmp_8_data_rsci_bcwt | tmp_8_data_rsci_biwt))
          | tmp_8_data_rsci_bdwt);
      tmp_8_data_rsci_douta_d_bfwt_15_0 <= tmp_8_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_8_data_rsci_oswt, tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_8_data_rsci_biwt,
      tmp_8_data_rsci_bdwt, tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_8_data_rsci_biwt_pff,
      tmp_8_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_8_data_rsci_oswt;
  input tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_8_data_rsci_biwt;
  output tmp_8_data_rsci_bdwt;
  output tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_8_data_rsci_biwt_pff;
  input tmp_8_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_8_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_8_data_rsci_bdwt = tmp_8_data_rsci_oswt & core_wen;
  assign tmp_8_data_rsci_biwt = (~ core_wten) & tmp_8_data_rsci_oswt;
  assign tmp_8_data_rsci_biwt_pff = tmp_8_data_rsci_tiswt0_pff;
  assign tmp_8_data_rsci_tiswt0_pff = core_wen & tmp_8_data_rsci_oswt_pff;
  assign tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_8_data_rsci_tiswt0_pff;
  assign tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_8_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_dp
    (
  clk, rst, tmp_7_data_rsci_addra_d, tmp_7_data_rsci_addrb_d, tmp_7_data_rsci_douta_d,
      tmp_7_data_rsci_addra_d_core, tmp_7_data_rsci_addrb_d_core, tmp_7_data_rsci_douta_d_mxwt,
      tmp_7_data_rsci_biwt, tmp_7_data_rsci_bdwt, tmp_7_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_7_data_rsci_addra_d;
  output [7:0] tmp_7_data_rsci_addrb_d;
  input [63:0] tmp_7_data_rsci_douta_d;
  input [7:0] tmp_7_data_rsci_addra_d_core;
  input [7:0] tmp_7_data_rsci_addrb_d_core;
  output [15:0] tmp_7_data_rsci_douta_d_mxwt;
  input tmp_7_data_rsci_biwt;
  input tmp_7_data_rsci_bdwt;
  input tmp_7_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_7_data_rsci_bcwt;
  reg [15:0] tmp_7_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_7_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_7_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_7_data_rsci_douta_d[15:0]),
      tmp_7_data_rsci_douta_d_bfwt_15_0, tmp_7_data_rsci_bcwt);
  assign tmp_7_data_rsci_douta_d_mxwt = tmp_7_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_7_data_rsci_addra_d = {(~ tmp_7_data_rsci_biwt_pff) , (tmp_7_data_rsci_addra_d_core[6:0])};
  assign tmp_7_data_rsci_addrb_d = {(~ tmp_7_data_rsci_biwt_pff) , (tmp_7_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_7_data_rsci_bcwt <= 1'b0;
      tmp_7_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_7_data_rsci_bcwt <= ~((~(tmp_7_data_rsci_bcwt | tmp_7_data_rsci_biwt))
          | tmp_7_data_rsci_bdwt);
      tmp_7_data_rsci_douta_d_bfwt_15_0 <= tmp_7_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_7_data_rsci_oswt, tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_7_data_rsci_biwt,
      tmp_7_data_rsci_bdwt, tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_7_data_rsci_biwt_pff,
      tmp_7_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_7_data_rsci_oswt;
  input tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_7_data_rsci_biwt;
  output tmp_7_data_rsci_bdwt;
  output tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_7_data_rsci_biwt_pff;
  input tmp_7_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_7_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_7_data_rsci_bdwt = tmp_7_data_rsci_oswt & core_wen;
  assign tmp_7_data_rsci_biwt = (~ core_wten) & tmp_7_data_rsci_oswt;
  assign tmp_7_data_rsci_biwt_pff = tmp_7_data_rsci_tiswt0_pff;
  assign tmp_7_data_rsci_tiswt0_pff = core_wen & tmp_7_data_rsci_oswt_pff;
  assign tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_7_data_rsci_tiswt0_pff;
  assign tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_7_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_dp
    (
  clk, rst, tmp_6_data_rsci_addra_d, tmp_6_data_rsci_addrb_d, tmp_6_data_rsci_douta_d,
      tmp_6_data_rsci_addra_d_core, tmp_6_data_rsci_addrb_d_core, tmp_6_data_rsci_douta_d_mxwt,
      tmp_6_data_rsci_biwt, tmp_6_data_rsci_bdwt, tmp_6_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_6_data_rsci_addra_d;
  output [7:0] tmp_6_data_rsci_addrb_d;
  input [63:0] tmp_6_data_rsci_douta_d;
  input [7:0] tmp_6_data_rsci_addra_d_core;
  input [7:0] tmp_6_data_rsci_addrb_d_core;
  output [15:0] tmp_6_data_rsci_douta_d_mxwt;
  input tmp_6_data_rsci_biwt;
  input tmp_6_data_rsci_bdwt;
  input tmp_6_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_6_data_rsci_bcwt;
  reg [15:0] tmp_6_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_6_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_6_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_6_data_rsci_douta_d[15:0]),
      tmp_6_data_rsci_douta_d_bfwt_15_0, tmp_6_data_rsci_bcwt);
  assign tmp_6_data_rsci_douta_d_mxwt = tmp_6_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_6_data_rsci_addra_d = {(~ tmp_6_data_rsci_biwt_pff) , (tmp_6_data_rsci_addra_d_core[6:0])};
  assign tmp_6_data_rsci_addrb_d = {(~ tmp_6_data_rsci_biwt_pff) , (tmp_6_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_6_data_rsci_bcwt <= 1'b0;
      tmp_6_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_6_data_rsci_bcwt <= ~((~(tmp_6_data_rsci_bcwt | tmp_6_data_rsci_biwt))
          | tmp_6_data_rsci_bdwt);
      tmp_6_data_rsci_douta_d_bfwt_15_0 <= tmp_6_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_6_data_rsci_oswt, tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_6_data_rsci_biwt,
      tmp_6_data_rsci_bdwt, tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_6_data_rsci_biwt_pff,
      tmp_6_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_6_data_rsci_oswt;
  input tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_6_data_rsci_biwt;
  output tmp_6_data_rsci_bdwt;
  output tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_6_data_rsci_biwt_pff;
  input tmp_6_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_6_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_6_data_rsci_bdwt = tmp_6_data_rsci_oswt & core_wen;
  assign tmp_6_data_rsci_biwt = (~ core_wten) & tmp_6_data_rsci_oswt;
  assign tmp_6_data_rsci_biwt_pff = tmp_6_data_rsci_tiswt0_pff;
  assign tmp_6_data_rsci_tiswt0_pff = core_wen & tmp_6_data_rsci_oswt_pff;
  assign tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_6_data_rsci_tiswt0_pff;
  assign tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_6_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_dp
    (
  clk, rst, tmp_5_data_rsci_addra_d, tmp_5_data_rsci_addrb_d, tmp_5_data_rsci_douta_d,
      tmp_5_data_rsci_addra_d_core, tmp_5_data_rsci_addrb_d_core, tmp_5_data_rsci_douta_d_mxwt,
      tmp_5_data_rsci_biwt, tmp_5_data_rsci_bdwt, tmp_5_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_5_data_rsci_addra_d;
  output [7:0] tmp_5_data_rsci_addrb_d;
  input [63:0] tmp_5_data_rsci_douta_d;
  input [7:0] tmp_5_data_rsci_addra_d_core;
  input [7:0] tmp_5_data_rsci_addrb_d_core;
  output [15:0] tmp_5_data_rsci_douta_d_mxwt;
  input tmp_5_data_rsci_biwt;
  input tmp_5_data_rsci_bdwt;
  input tmp_5_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_5_data_rsci_bcwt;
  reg [15:0] tmp_5_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_5_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_5_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_5_data_rsci_douta_d[15:0]),
      tmp_5_data_rsci_douta_d_bfwt_15_0, tmp_5_data_rsci_bcwt);
  assign tmp_5_data_rsci_douta_d_mxwt = tmp_5_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_5_data_rsci_addra_d = {(~ tmp_5_data_rsci_biwt_pff) , (tmp_5_data_rsci_addra_d_core[6:0])};
  assign tmp_5_data_rsci_addrb_d = {(~ tmp_5_data_rsci_biwt_pff) , (tmp_5_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_5_data_rsci_bcwt <= 1'b0;
      tmp_5_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_5_data_rsci_bcwt <= ~((~(tmp_5_data_rsci_bcwt | tmp_5_data_rsci_biwt))
          | tmp_5_data_rsci_bdwt);
      tmp_5_data_rsci_douta_d_bfwt_15_0 <= tmp_5_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_5_data_rsci_oswt, tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_5_data_rsci_biwt,
      tmp_5_data_rsci_bdwt, tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_5_data_rsci_biwt_pff,
      tmp_5_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_5_data_rsci_oswt;
  input tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_5_data_rsci_biwt;
  output tmp_5_data_rsci_bdwt;
  output tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_5_data_rsci_biwt_pff;
  input tmp_5_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_5_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_5_data_rsci_bdwt = tmp_5_data_rsci_oswt & core_wen;
  assign tmp_5_data_rsci_biwt = (~ core_wten) & tmp_5_data_rsci_oswt;
  assign tmp_5_data_rsci_biwt_pff = tmp_5_data_rsci_tiswt0_pff;
  assign tmp_5_data_rsci_tiswt0_pff = core_wen & tmp_5_data_rsci_oswt_pff;
  assign tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_5_data_rsci_tiswt0_pff;
  assign tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_5_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_dp
    (
  clk, rst, tmp_4_data_rsci_addra_d, tmp_4_data_rsci_addrb_d, tmp_4_data_rsci_douta_d,
      tmp_4_data_rsci_addra_d_core, tmp_4_data_rsci_addrb_d_core, tmp_4_data_rsci_douta_d_mxwt,
      tmp_4_data_rsci_biwt, tmp_4_data_rsci_bdwt, tmp_4_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_4_data_rsci_addra_d;
  output [7:0] tmp_4_data_rsci_addrb_d;
  input [63:0] tmp_4_data_rsci_douta_d;
  input [7:0] tmp_4_data_rsci_addra_d_core;
  input [7:0] tmp_4_data_rsci_addrb_d_core;
  output [15:0] tmp_4_data_rsci_douta_d_mxwt;
  input tmp_4_data_rsci_biwt;
  input tmp_4_data_rsci_bdwt;
  input tmp_4_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_4_data_rsci_bcwt;
  reg [15:0] tmp_4_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_4_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_4_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_4_data_rsci_douta_d[15:0]),
      tmp_4_data_rsci_douta_d_bfwt_15_0, tmp_4_data_rsci_bcwt);
  assign tmp_4_data_rsci_douta_d_mxwt = tmp_4_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_4_data_rsci_addra_d = {(~ tmp_4_data_rsci_biwt_pff) , (tmp_4_data_rsci_addra_d_core[6:0])};
  assign tmp_4_data_rsci_addrb_d = {(~ tmp_4_data_rsci_biwt_pff) , (tmp_4_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_4_data_rsci_bcwt <= 1'b0;
      tmp_4_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_4_data_rsci_bcwt <= ~((~(tmp_4_data_rsci_bcwt | tmp_4_data_rsci_biwt))
          | tmp_4_data_rsci_bdwt);
      tmp_4_data_rsci_douta_d_bfwt_15_0 <= tmp_4_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_4_data_rsci_oswt, tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_4_data_rsci_biwt,
      tmp_4_data_rsci_bdwt, tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_4_data_rsci_biwt_pff,
      tmp_4_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_4_data_rsci_oswt;
  input tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_4_data_rsci_biwt;
  output tmp_4_data_rsci_bdwt;
  output tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_4_data_rsci_biwt_pff;
  input tmp_4_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_4_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_4_data_rsci_bdwt = tmp_4_data_rsci_oswt & core_wen;
  assign tmp_4_data_rsci_biwt = (~ core_wten) & tmp_4_data_rsci_oswt;
  assign tmp_4_data_rsci_biwt_pff = tmp_4_data_rsci_tiswt0_pff;
  assign tmp_4_data_rsci_tiswt0_pff = core_wen & tmp_4_data_rsci_oswt_pff;
  assign tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_4_data_rsci_tiswt0_pff;
  assign tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_4_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_dp
    (
  clk, rst, tmp_3_data_rsci_addra_d, tmp_3_data_rsci_addrb_d, tmp_3_data_rsci_douta_d,
      tmp_3_data_rsci_addra_d_core, tmp_3_data_rsci_addrb_d_core, tmp_3_data_rsci_douta_d_mxwt,
      tmp_3_data_rsci_biwt, tmp_3_data_rsci_bdwt, tmp_3_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_3_data_rsci_addra_d;
  output [7:0] tmp_3_data_rsci_addrb_d;
  input [63:0] tmp_3_data_rsci_douta_d;
  input [7:0] tmp_3_data_rsci_addra_d_core;
  input [7:0] tmp_3_data_rsci_addrb_d_core;
  output [15:0] tmp_3_data_rsci_douta_d_mxwt;
  input tmp_3_data_rsci_biwt;
  input tmp_3_data_rsci_bdwt;
  input tmp_3_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_3_data_rsci_bcwt;
  reg [15:0] tmp_3_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_3_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_3_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_3_data_rsci_douta_d[15:0]),
      tmp_3_data_rsci_douta_d_bfwt_15_0, tmp_3_data_rsci_bcwt);
  assign tmp_3_data_rsci_douta_d_mxwt = tmp_3_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_3_data_rsci_addra_d = {(~ tmp_3_data_rsci_biwt_pff) , (tmp_3_data_rsci_addra_d_core[6:0])};
  assign tmp_3_data_rsci_addrb_d = {(~ tmp_3_data_rsci_biwt_pff) , (tmp_3_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_3_data_rsci_bcwt <= 1'b0;
      tmp_3_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_3_data_rsci_bcwt <= ~((~(tmp_3_data_rsci_bcwt | tmp_3_data_rsci_biwt))
          | tmp_3_data_rsci_bdwt);
      tmp_3_data_rsci_douta_d_bfwt_15_0 <= tmp_3_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_3_data_rsci_oswt, tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_3_data_rsci_biwt,
      tmp_3_data_rsci_bdwt, tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_3_data_rsci_biwt_pff,
      tmp_3_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_3_data_rsci_oswt;
  input tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_3_data_rsci_biwt;
  output tmp_3_data_rsci_bdwt;
  output tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_3_data_rsci_biwt_pff;
  input tmp_3_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_3_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_3_data_rsci_bdwt = tmp_3_data_rsci_oswt & core_wen;
  assign tmp_3_data_rsci_biwt = (~ core_wten) & tmp_3_data_rsci_oswt;
  assign tmp_3_data_rsci_biwt_pff = tmp_3_data_rsci_tiswt0_pff;
  assign tmp_3_data_rsci_tiswt0_pff = core_wen & tmp_3_data_rsci_oswt_pff;
  assign tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_3_data_rsci_tiswt0_pff;
  assign tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_3_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_dp
    (
  clk, rst, tmp_2_data_rsci_addra_d, tmp_2_data_rsci_addrb_d, tmp_2_data_rsci_douta_d,
      tmp_2_data_rsci_addra_d_core, tmp_2_data_rsci_addrb_d_core, tmp_2_data_rsci_douta_d_mxwt,
      tmp_2_data_rsci_biwt, tmp_2_data_rsci_bdwt, tmp_2_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_2_data_rsci_addra_d;
  output [7:0] tmp_2_data_rsci_addrb_d;
  input [63:0] tmp_2_data_rsci_douta_d;
  input [7:0] tmp_2_data_rsci_addra_d_core;
  input [7:0] tmp_2_data_rsci_addrb_d_core;
  output [15:0] tmp_2_data_rsci_douta_d_mxwt;
  input tmp_2_data_rsci_biwt;
  input tmp_2_data_rsci_bdwt;
  input tmp_2_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_2_data_rsci_bcwt;
  reg [15:0] tmp_2_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_2_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_2_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_2_data_rsci_douta_d[15:0]),
      tmp_2_data_rsci_douta_d_bfwt_15_0, tmp_2_data_rsci_bcwt);
  assign tmp_2_data_rsci_douta_d_mxwt = tmp_2_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_2_data_rsci_addra_d = {(~ tmp_2_data_rsci_biwt_pff) , (tmp_2_data_rsci_addra_d_core[6:0])};
  assign tmp_2_data_rsci_addrb_d = {(~ tmp_2_data_rsci_biwt_pff) , (tmp_2_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_2_data_rsci_bcwt <= 1'b0;
      tmp_2_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_2_data_rsci_bcwt <= ~((~(tmp_2_data_rsci_bcwt | tmp_2_data_rsci_biwt))
          | tmp_2_data_rsci_bdwt);
      tmp_2_data_rsci_douta_d_bfwt_15_0 <= tmp_2_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_2_data_rsci_oswt, tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_2_data_rsci_biwt,
      tmp_2_data_rsci_bdwt, tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_2_data_rsci_biwt_pff,
      tmp_2_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_2_data_rsci_oswt;
  input tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_2_data_rsci_biwt;
  output tmp_2_data_rsci_bdwt;
  output tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_2_data_rsci_biwt_pff;
  input tmp_2_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_2_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_2_data_rsci_bdwt = tmp_2_data_rsci_oswt & core_wen;
  assign tmp_2_data_rsci_biwt = (~ core_wten) & tmp_2_data_rsci_oswt;
  assign tmp_2_data_rsci_biwt_pff = tmp_2_data_rsci_tiswt0_pff;
  assign tmp_2_data_rsci_tiswt0_pff = core_wen & tmp_2_data_rsci_oswt_pff;
  assign tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_2_data_rsci_tiswt0_pff;
  assign tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_2_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_dp
    (
  clk, rst, tmp_1_data_rsci_addra_d, tmp_1_data_rsci_addrb_d, tmp_1_data_rsci_douta_d,
      tmp_1_data_rsci_addra_d_core, tmp_1_data_rsci_addrb_d_core, tmp_1_data_rsci_douta_d_mxwt,
      tmp_1_data_rsci_biwt, tmp_1_data_rsci_bdwt, tmp_1_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_1_data_rsci_addra_d;
  output [7:0] tmp_1_data_rsci_addrb_d;
  input [63:0] tmp_1_data_rsci_douta_d;
  input [7:0] tmp_1_data_rsci_addra_d_core;
  input [7:0] tmp_1_data_rsci_addrb_d_core;
  output [15:0] tmp_1_data_rsci_douta_d_mxwt;
  input tmp_1_data_rsci_biwt;
  input tmp_1_data_rsci_bdwt;
  input tmp_1_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_1_data_rsci_bcwt;
  reg [15:0] tmp_1_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_1_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_1_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_1_data_rsci_douta_d[15:0]),
      tmp_1_data_rsci_douta_d_bfwt_15_0, tmp_1_data_rsci_bcwt);
  assign tmp_1_data_rsci_douta_d_mxwt = tmp_1_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_1_data_rsci_addra_d = {(~ tmp_1_data_rsci_biwt_pff) , (tmp_1_data_rsci_addra_d_core[6:0])};
  assign tmp_1_data_rsci_addrb_d = {(~ tmp_1_data_rsci_biwt_pff) , (tmp_1_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_1_data_rsci_bcwt <= 1'b0;
      tmp_1_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_1_data_rsci_bcwt <= ~((~(tmp_1_data_rsci_bcwt | tmp_1_data_rsci_biwt))
          | tmp_1_data_rsci_bdwt);
      tmp_1_data_rsci_douta_d_bfwt_15_0 <= tmp_1_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_1_data_rsci_oswt, tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_1_data_rsci_biwt,
      tmp_1_data_rsci_bdwt, tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_1_data_rsci_biwt_pff,
      tmp_1_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_1_data_rsci_oswt;
  input tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_1_data_rsci_biwt;
  output tmp_1_data_rsci_bdwt;
  output tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_1_data_rsci_biwt_pff;
  input tmp_1_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_1_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_1_data_rsci_bdwt = tmp_1_data_rsci_oswt & core_wen;
  assign tmp_1_data_rsci_biwt = (~ core_wten) & tmp_1_data_rsci_oswt;
  assign tmp_1_data_rsci_biwt_pff = tmp_1_data_rsci_tiswt0_pff;
  assign tmp_1_data_rsci_tiswt0_pff = core_wen & tmp_1_data_rsci_oswt_pff;
  assign tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_1_data_rsci_tiswt0_pff;
  assign tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_1_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_dp
    (
  clk, rst, tmp_0_data_rsci_addra_d, tmp_0_data_rsci_addrb_d, tmp_0_data_rsci_douta_d,
      tmp_0_data_rsci_addra_d_core, tmp_0_data_rsci_addrb_d_core, tmp_0_data_rsci_douta_d_mxwt,
      tmp_0_data_rsci_biwt, tmp_0_data_rsci_bdwt, tmp_0_data_rsci_biwt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_0_data_rsci_addra_d;
  output [7:0] tmp_0_data_rsci_addrb_d;
  input [63:0] tmp_0_data_rsci_douta_d;
  input [7:0] tmp_0_data_rsci_addra_d_core;
  input [7:0] tmp_0_data_rsci_addrb_d_core;
  output [15:0] tmp_0_data_rsci_douta_d_mxwt;
  input tmp_0_data_rsci_biwt;
  input tmp_0_data_rsci_bdwt;
  input tmp_0_data_rsci_biwt_pff;


  // Interconnect Declarations
  reg tmp_0_data_rsci_bcwt;
  reg [15:0] tmp_0_data_rsci_douta_d_bfwt_15_0;
  wire [15:0] tmp_0_data_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_0_data_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((tmp_0_data_rsci_douta_d[15:0]),
      tmp_0_data_rsci_douta_d_bfwt_15_0, tmp_0_data_rsci_bcwt);
  assign tmp_0_data_rsci_douta_d_mxwt = tmp_0_data_rsci_douta_d_mxwt_opt_15_0;
  assign tmp_0_data_rsci_addra_d = {(~ tmp_0_data_rsci_biwt_pff) , (tmp_0_data_rsci_addra_d_core[6:0])};
  assign tmp_0_data_rsci_addrb_d = {(~ tmp_0_data_rsci_biwt_pff) , (tmp_0_data_rsci_addrb_d_core[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_0_data_rsci_bcwt <= 1'b0;
      tmp_0_data_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      tmp_0_data_rsci_bcwt <= ~((~(tmp_0_data_rsci_bcwt | tmp_0_data_rsci_biwt))
          | tmp_0_data_rsci_bdwt);
      tmp_0_data_rsci_douta_d_bfwt_15_0 <= tmp_0_data_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_ctrl
    (
  core_wen, core_wten, tmp_0_data_rsci_oswt, tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_0_data_rsci_biwt,
      tmp_0_data_rsci_bdwt, tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct,
      tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct, tmp_0_data_rsci_biwt_pff,
      tmp_0_data_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input tmp_0_data_rsci_oswt;
  input tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  output tmp_0_data_rsci_biwt;
  output tmp_0_data_rsci_bdwt;
  output tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  output tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  output tmp_0_data_rsci_biwt_pff;
  input tmp_0_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_0_data_rsci_tiswt0_pff;


  // Interconnect Declarations for Component Instantiations 
  assign tmp_0_data_rsci_bdwt = tmp_0_data_rsci_oswt & core_wen;
  assign tmp_0_data_rsci_biwt = (~ core_wten) & tmp_0_data_rsci_oswt;
  assign tmp_0_data_rsci_biwt_pff = tmp_0_data_rsci_tiswt0_pff;
  assign tmp_0_data_rsci_tiswt0_pff = core_wen & tmp_0_data_rsci_oswt_pff;
  assign tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct = tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      & tmp_0_data_rsci_tiswt0_pff;
  assign tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      & tmp_0_data_rsci_tiswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_dout_17_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_dout_17_rsc_wait_ctrl
    (
  dout_17_rsci_dinb_d_core_sct_pff, dout_17_rsci_iswt0_pff, core_wten_pff
);
  output dout_17_rsci_dinb_d_core_sct_pff;
  input dout_17_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_17_rsci_dinb_d_core_sct_pff = dout_17_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_dout_16_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_dout_16_rsc_wait_ctrl
    (
  dout_16_rsci_dinb_d_core_sct_pff, dout_16_rsci_iswt0_pff, core_wten_pff
);
  output dout_16_rsci_dinb_d_core_sct_pff;
  input dout_16_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_16_rsci_dinb_d_core_sct_pff = dout_16_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_dout_15_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_dout_15_rsc_wait_ctrl
    (
  dout_15_rsci_dinb_d_core_sct_pff, dout_15_rsci_iswt0_pff, core_wten_pff
);
  output dout_15_rsci_dinb_d_core_sct_pff;
  input dout_15_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_15_rsci_dinb_d_core_sct_pff = dout_15_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_dout_14_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_dout_14_rsc_wait_ctrl
    (
  dout_14_rsci_dinb_d_core_sct_pff, dout_14_rsci_iswt0_pff, core_wten_pff
);
  output dout_14_rsci_dinb_d_core_sct_pff;
  input dout_14_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_14_rsci_dinb_d_core_sct_pff = dout_14_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_dout_13_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_dout_13_rsc_wait_ctrl
    (
  dout_13_rsci_dinb_d_core_sct_pff, dout_13_rsci_iswt0_pff, core_wten_pff
);
  output dout_13_rsci_dinb_d_core_sct_pff;
  input dout_13_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_13_rsci_dinb_d_core_sct_pff = dout_13_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_dout_12_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_dout_12_rsc_wait_ctrl
    (
  dout_12_rsci_dinb_d_core_sct_pff, dout_12_rsci_iswt0_pff, core_wten_pff
);
  output dout_12_rsci_dinb_d_core_sct_pff;
  input dout_12_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_12_rsci_dinb_d_core_sct_pff = dout_12_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_dout_11_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_dout_11_rsc_wait_ctrl
    (
  dout_11_rsci_dinb_d_core_sct_pff, dout_11_rsci_iswt0_pff, core_wten_pff
);
  output dout_11_rsci_dinb_d_core_sct_pff;
  input dout_11_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_11_rsci_dinb_d_core_sct_pff = dout_11_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_dout_10_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_dout_10_rsc_wait_ctrl
    (
  dout_10_rsci_dinb_d_core_sct_pff, dout_10_rsci_iswt0_pff, core_wten_pff
);
  output dout_10_rsci_dinb_d_core_sct_pff;
  input dout_10_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_10_rsci_dinb_d_core_sct_pff = dout_10_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_dout_9_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_dout_9_rsc_wait_ctrl
    (
  dout_9_rsci_dinb_d_core_sct_pff, dout_9_rsci_iswt0_pff, core_wten_pff
);
  output dout_9_rsci_dinb_d_core_sct_pff;
  input dout_9_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_9_rsci_dinb_d_core_sct_pff = dout_9_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_dout_8_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_dout_8_rsc_wait_ctrl
    (
  dout_8_rsci_dinb_d_core_sct_pff, dout_8_rsci_iswt0_pff, core_wten_pff
);
  output dout_8_rsci_dinb_d_core_sct_pff;
  input dout_8_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_8_rsci_dinb_d_core_sct_pff = dout_8_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_dout_7_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_dout_7_rsc_wait_ctrl
    (
  dout_7_rsci_dinb_d_core_sct_pff, dout_7_rsci_iswt0_pff, core_wten_pff
);
  output dout_7_rsci_dinb_d_core_sct_pff;
  input dout_7_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_7_rsci_dinb_d_core_sct_pff = dout_7_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_dout_6_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_dout_6_rsc_wait_ctrl
    (
  dout_6_rsci_dinb_d_core_sct_pff, dout_6_rsci_iswt0_pff, core_wten_pff
);
  output dout_6_rsci_dinb_d_core_sct_pff;
  input dout_6_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_6_rsci_dinb_d_core_sct_pff = dout_6_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_dout_5_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_dout_5_rsc_wait_ctrl
    (
  dout_5_rsci_dinb_d_core_sct_pff, dout_5_rsci_iswt0_pff, core_wten_pff
);
  output dout_5_rsci_dinb_d_core_sct_pff;
  input dout_5_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_5_rsci_dinb_d_core_sct_pff = dout_5_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_dout_4_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_dout_4_rsc_wait_ctrl
    (
  dout_4_rsci_dinb_d_core_sct_pff, dout_4_rsci_iswt0_pff, core_wten_pff
);
  output dout_4_rsci_dinb_d_core_sct_pff;
  input dout_4_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_4_rsci_dinb_d_core_sct_pff = dout_4_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_dout_3_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_dout_3_rsc_wait_ctrl
    (
  dout_3_rsci_dinb_d_core_sct_pff, dout_3_rsci_iswt0_pff, core_wten_pff
);
  output dout_3_rsci_dinb_d_core_sct_pff;
  input dout_3_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_3_rsci_dinb_d_core_sct_pff = dout_3_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_dout_2_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_dout_2_rsc_wait_ctrl
    (
  dout_2_rsci_dinb_d_core_sct_pff, dout_2_rsci_iswt0_pff, core_wten_pff
);
  output dout_2_rsci_dinb_d_core_sct_pff;
  input dout_2_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_2_rsci_dinb_d_core_sct_pff = dout_2_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_dout_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_dout_1_rsc_wait_ctrl
    (
  dout_1_rsci_dinb_d_core_sct_pff, dout_1_rsci_iswt0_pff, core_wten_pff
);
  output dout_1_rsci_dinb_d_core_sct_pff;
  input dout_1_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_1_rsci_dinb_d_core_sct_pff = dout_1_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_dout_0_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_dout_0_rsc_wait_ctrl
    (
  dout_0_rsci_dinb_d_core_sct_pff, dout_0_rsci_iswt0_pff, core_wten_pff
);
  output dout_0_rsci_dinb_d_core_sct_pff;
  input dout_0_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_0_rsci_dinb_d_core_sct_pff = dout_0_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci_din_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci_din_wait_dp (
  clk, rst, din_rsci_oswt, din_rsci_wen_comp, din_rsci_d_mxwt, din_rsci_biwt, din_rsci_bdwt,
      din_rsci_d
);
  input clk;
  input rst;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [15:0] din_rsci_d_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  input [15:0] din_rsci_d;


  // Interconnect Declarations
  reg din_rsci_bcwt;
  reg [15:0] din_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_wen_comp = (~ din_rsci_oswt) | din_rsci_biwt | din_rsci_bcwt;
  assign din_rsci_d_mxwt = MUX_v_16_2_2(din_rsci_d, din_rsci_d_bfwt, din_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsci_bcwt <= 1'b0;
      din_rsci_d_bfwt <= 16'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
      din_rsci_d_bfwt <= din_rsci_d_mxwt;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci_din_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci_din_wait_ctrl (
  clk, rst, core_wen, din_rsci_oswt, core_wten, din_rsci_biwt, din_rsci_bdwt, din_rsci_ld_core_sct,
      din_rsci_vd
);
  input clk;
  input rst;
  input core_wen;
  input din_rsci_oswt;
  input core_wten;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  output din_rsci_ld_core_sct;
  input din_rsci_vd;


  // Interconnect Declarations
  wire din_rsci_ogwt;
  wire din_rsci_pdswt0;
  reg din_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_pdswt0 = (~ core_wten) & din_rsci_oswt;
  assign din_rsci_biwt = din_rsci_ogwt & din_rsci_vd;
  assign din_rsci_ogwt = din_rsci_pdswt0 | din_rsci_icwt;
  assign din_rsci_bdwt = din_rsci_oswt & core_wen;
  assign din_rsci_ld_core_sct = din_rsci_oswt & din_rsci_ogwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsci_icwt <= 1'b0;
    end
    else begin
      din_rsci_icwt <= ~((~(din_rsci_icwt | din_rsci_pdswt0)) | din_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_55_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_55_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_17_and_nl;
  wire din_17_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_17_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_17_and_nl);
  assign din_17_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_17_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_54_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_54_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_16_and_nl;
  wire din_16_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_16_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_16_and_nl);
  assign din_16_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_16_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_53_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_53_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_15_and_nl;
  wire din_15_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_15_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_15_and_nl);
  assign din_15_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_15_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_52_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_52_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_14_and_nl;
  wire din_14_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_14_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_14_and_nl);
  assign din_14_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_14_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_51_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_51_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_13_and_nl;
  wire din_13_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_13_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_13_and_nl);
  assign din_13_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_13_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_50_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_50_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_12_and_nl;
  wire din_12_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_12_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_12_and_nl);
  assign din_12_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_12_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_49_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_49_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_11_and_nl;
  wire din_11_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_11_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_11_and_nl);
  assign din_11_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_11_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_48_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_48_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_10_and_nl;
  wire din_10_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_10_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_10_and_nl);
  assign din_10_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_10_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_47_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_47_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_9_and_nl;
  wire din_9_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_9_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_9_and_nl);
  assign din_9_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_9_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_46_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_46_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_8_and_nl;
  wire din_8_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_8_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_8_and_nl);
  assign din_8_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_8_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_45_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_45_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_7_and_nl;
  wire din_7_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_7_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_7_and_nl);
  assign din_7_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_7_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_44_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_44_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_6_and_nl;
  wire din_6_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_6_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_6_and_nl);
  assign din_6_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_6_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_43_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_43_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_5_and_nl;
  wire din_5_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_5_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_5_and_nl);
  assign din_5_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_5_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_42_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_42_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_4_and_nl;
  wire din_4_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_4_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_4_and_nl);
  assign din_4_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_4_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_41_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_41_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_3_and_nl;
  wire din_3_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_3_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_3_and_nl);
  assign din_3_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_3_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_40_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_40_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_2_and_nl;
  wire din_2_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_2_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_2_and_nl);
  assign din_2_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_2_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_39_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_39_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_1_and_nl;
  wire din_1_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_1_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_1_and_nl);
  assign din_1_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_1_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_38_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_38_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_0_and_nl;
  wire din_0_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_0_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_0_and_nl);
  assign din_0_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_0_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_staller
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_staller (
  clk, rst, core_wen, core_wten, dout_rsci_wen_comp, din_17_rsc_req_obj_wen_comp,
      din_16_rsc_req_obj_wen_comp, din_15_rsc_req_obj_wen_comp, din_14_rsc_req_obj_wen_comp,
      din_13_rsc_req_obj_wen_comp, din_12_rsc_req_obj_wen_comp, din_11_rsc_req_obj_wen_comp,
      din_10_rsc_req_obj_wen_comp, din_9_rsc_req_obj_wen_comp, din_8_rsc_req_obj_wen_comp,
      din_7_rsc_req_obj_wen_comp, din_6_rsc_req_obj_wen_comp, din_5_rsc_req_obj_wen_comp,
      din_4_rsc_req_obj_wen_comp, din_3_rsc_req_obj_wen_comp, din_2_rsc_req_obj_wen_comp,
      din_1_rsc_req_obj_wen_comp, din_0_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input dout_rsci_wen_comp;
  input din_17_rsc_req_obj_wen_comp;
  input din_16_rsc_req_obj_wen_comp;
  input din_15_rsc_req_obj_wen_comp;
  input din_14_rsc_req_obj_wen_comp;
  input din_13_rsc_req_obj_wen_comp;
  input din_12_rsc_req_obj_wen_comp;
  input din_11_rsc_req_obj_wen_comp;
  input din_10_rsc_req_obj_wen_comp;
  input din_9_rsc_req_obj_wen_comp;
  input din_8_rsc_req_obj_wen_comp;
  input din_7_rsc_req_obj_wen_comp;
  input din_6_rsc_req_obj_wen_comp;
  input din_5_rsc_req_obj_wen_comp;
  input din_4_rsc_req_obj_wen_comp;
  input din_3_rsc_req_obj_wen_comp;
  input din_2_rsc_req_obj_wen_comp;
  input din_1_rsc_req_obj_wen_comp;
  input din_0_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = dout_rsci_wen_comp & din_17_rsc_req_obj_wen_comp & din_16_rsc_req_obj_wen_comp
      & din_15_rsc_req_obj_wen_comp & din_14_rsc_req_obj_wen_comp & din_13_rsc_req_obj_wen_comp
      & din_12_rsc_req_obj_wen_comp & din_11_rsc_req_obj_wen_comp & din_10_rsc_req_obj_wen_comp
      & din_9_rsc_req_obj_wen_comp & din_8_rsc_req_obj_wen_comp & din_7_rsc_req_obj_wen_comp
      & din_6_rsc_req_obj_wen_comp & din_5_rsc_req_obj_wen_comp & din_4_rsc_req_obj_wen_comp
      & din_3_rsc_req_obj_wen_comp & din_2_rsc_req_obj_wen_comp & din_1_rsc_req_obj_wen_comp
      & din_0_rsc_req_obj_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj_din_0_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj_din_0_rsc_req_wait_dp
    (
  clk, rst, din_0_rsc_req_obj_oswt, din_0_rsc_req_obj_wen_comp, din_0_rsc_req_obj_biwt,
      din_0_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_0_rsc_req_obj_oswt;
  output din_0_rsc_req_obj_wen_comp;
  input din_0_rsc_req_obj_biwt;
  input din_0_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_0_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_0_rsc_req_obj_wen_comp = (~ din_0_rsc_req_obj_oswt) | din_0_rsc_req_obj_biwt
      | din_0_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_0_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_0_rsc_req_obj_bcwt <= ~((~(din_0_rsc_req_obj_bcwt | din_0_rsc_req_obj_biwt))
          | din_0_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj_din_0_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj_din_0_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_0_rsc_req_obj_oswt, din_0_rsc_req_obj_vd, din_0_rsc_req_obj_biwt,
      din_0_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_0_rsc_req_obj_oswt;
  input din_0_rsc_req_obj_vd;
  output din_0_rsc_req_obj_biwt;
  output din_0_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_0_rsc_req_obj_pdswt0;
  reg din_0_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_0_rsc_req_obj_pdswt0 = (~ core_wten) & din_0_rsc_req_obj_oswt;
  assign din_0_rsc_req_obj_biwt = (din_0_rsc_req_obj_pdswt0 | din_0_rsc_req_obj_icwt)
      & din_0_rsc_req_obj_vd;
  assign din_0_rsc_req_obj_bdwt = din_0_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_0_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_0_rsc_req_obj_icwt <= ~((~(din_0_rsc_req_obj_icwt | din_0_rsc_req_obj_pdswt0))
          | din_0_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj_din_1_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj_din_1_rsc_req_wait_dp
    (
  clk, rst, din_1_rsc_req_obj_oswt, din_1_rsc_req_obj_wen_comp, din_1_rsc_req_obj_biwt,
      din_1_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_1_rsc_req_obj_oswt;
  output din_1_rsc_req_obj_wen_comp;
  input din_1_rsc_req_obj_biwt;
  input din_1_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_1_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_1_rsc_req_obj_wen_comp = (~ din_1_rsc_req_obj_oswt) | din_1_rsc_req_obj_biwt
      | din_1_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_1_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_1_rsc_req_obj_bcwt <= ~((~(din_1_rsc_req_obj_bcwt | din_1_rsc_req_obj_biwt))
          | din_1_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj_din_1_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj_din_1_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_1_rsc_req_obj_oswt, din_1_rsc_req_obj_vd, din_1_rsc_req_obj_biwt,
      din_1_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_1_rsc_req_obj_oswt;
  input din_1_rsc_req_obj_vd;
  output din_1_rsc_req_obj_biwt;
  output din_1_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_1_rsc_req_obj_pdswt0;
  reg din_1_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_1_rsc_req_obj_pdswt0 = (~ core_wten) & din_1_rsc_req_obj_oswt;
  assign din_1_rsc_req_obj_biwt = (din_1_rsc_req_obj_pdswt0 | din_1_rsc_req_obj_icwt)
      & din_1_rsc_req_obj_vd;
  assign din_1_rsc_req_obj_bdwt = din_1_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_1_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_1_rsc_req_obj_icwt <= ~((~(din_1_rsc_req_obj_icwt | din_1_rsc_req_obj_pdswt0))
          | din_1_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj_din_2_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj_din_2_rsc_req_wait_dp
    (
  clk, rst, din_2_rsc_req_obj_oswt, din_2_rsc_req_obj_wen_comp, din_2_rsc_req_obj_biwt,
      din_2_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_2_rsc_req_obj_oswt;
  output din_2_rsc_req_obj_wen_comp;
  input din_2_rsc_req_obj_biwt;
  input din_2_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_2_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_2_rsc_req_obj_wen_comp = (~ din_2_rsc_req_obj_oswt) | din_2_rsc_req_obj_biwt
      | din_2_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_2_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_2_rsc_req_obj_bcwt <= ~((~(din_2_rsc_req_obj_bcwt | din_2_rsc_req_obj_biwt))
          | din_2_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj_din_2_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj_din_2_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_2_rsc_req_obj_oswt, din_2_rsc_req_obj_vd, din_2_rsc_req_obj_biwt,
      din_2_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_2_rsc_req_obj_oswt;
  input din_2_rsc_req_obj_vd;
  output din_2_rsc_req_obj_biwt;
  output din_2_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_2_rsc_req_obj_pdswt0;
  reg din_2_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_2_rsc_req_obj_pdswt0 = (~ core_wten) & din_2_rsc_req_obj_oswt;
  assign din_2_rsc_req_obj_biwt = (din_2_rsc_req_obj_pdswt0 | din_2_rsc_req_obj_icwt)
      & din_2_rsc_req_obj_vd;
  assign din_2_rsc_req_obj_bdwt = din_2_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_2_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_2_rsc_req_obj_icwt <= ~((~(din_2_rsc_req_obj_icwt | din_2_rsc_req_obj_pdswt0))
          | din_2_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj_din_3_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj_din_3_rsc_req_wait_dp
    (
  clk, rst, din_3_rsc_req_obj_oswt, din_3_rsc_req_obj_wen_comp, din_3_rsc_req_obj_biwt,
      din_3_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_3_rsc_req_obj_oswt;
  output din_3_rsc_req_obj_wen_comp;
  input din_3_rsc_req_obj_biwt;
  input din_3_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_3_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_3_rsc_req_obj_wen_comp = (~ din_3_rsc_req_obj_oswt) | din_3_rsc_req_obj_biwt
      | din_3_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_3_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_3_rsc_req_obj_bcwt <= ~((~(din_3_rsc_req_obj_bcwt | din_3_rsc_req_obj_biwt))
          | din_3_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj_din_3_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj_din_3_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_3_rsc_req_obj_oswt, din_3_rsc_req_obj_vd, din_3_rsc_req_obj_biwt,
      din_3_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_3_rsc_req_obj_oswt;
  input din_3_rsc_req_obj_vd;
  output din_3_rsc_req_obj_biwt;
  output din_3_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_3_rsc_req_obj_pdswt0;
  reg din_3_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_3_rsc_req_obj_pdswt0 = (~ core_wten) & din_3_rsc_req_obj_oswt;
  assign din_3_rsc_req_obj_biwt = (din_3_rsc_req_obj_pdswt0 | din_3_rsc_req_obj_icwt)
      & din_3_rsc_req_obj_vd;
  assign din_3_rsc_req_obj_bdwt = din_3_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_3_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_3_rsc_req_obj_icwt <= ~((~(din_3_rsc_req_obj_icwt | din_3_rsc_req_obj_pdswt0))
          | din_3_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj_din_4_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj_din_4_rsc_req_wait_dp
    (
  clk, rst, din_4_rsc_req_obj_oswt, din_4_rsc_req_obj_wen_comp, din_4_rsc_req_obj_biwt,
      din_4_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_4_rsc_req_obj_oswt;
  output din_4_rsc_req_obj_wen_comp;
  input din_4_rsc_req_obj_biwt;
  input din_4_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_4_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_4_rsc_req_obj_wen_comp = (~ din_4_rsc_req_obj_oswt) | din_4_rsc_req_obj_biwt
      | din_4_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_4_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_4_rsc_req_obj_bcwt <= ~((~(din_4_rsc_req_obj_bcwt | din_4_rsc_req_obj_biwt))
          | din_4_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj_din_4_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj_din_4_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_4_rsc_req_obj_oswt, din_4_rsc_req_obj_vd, din_4_rsc_req_obj_biwt,
      din_4_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_4_rsc_req_obj_oswt;
  input din_4_rsc_req_obj_vd;
  output din_4_rsc_req_obj_biwt;
  output din_4_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_4_rsc_req_obj_pdswt0;
  reg din_4_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_4_rsc_req_obj_pdswt0 = (~ core_wten) & din_4_rsc_req_obj_oswt;
  assign din_4_rsc_req_obj_biwt = (din_4_rsc_req_obj_pdswt0 | din_4_rsc_req_obj_icwt)
      & din_4_rsc_req_obj_vd;
  assign din_4_rsc_req_obj_bdwt = din_4_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_4_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_4_rsc_req_obj_icwt <= ~((~(din_4_rsc_req_obj_icwt | din_4_rsc_req_obj_pdswt0))
          | din_4_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj_din_5_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj_din_5_rsc_req_wait_dp
    (
  clk, rst, din_5_rsc_req_obj_oswt, din_5_rsc_req_obj_wen_comp, din_5_rsc_req_obj_biwt,
      din_5_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_5_rsc_req_obj_oswt;
  output din_5_rsc_req_obj_wen_comp;
  input din_5_rsc_req_obj_biwt;
  input din_5_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_5_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_5_rsc_req_obj_wen_comp = (~ din_5_rsc_req_obj_oswt) | din_5_rsc_req_obj_biwt
      | din_5_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_5_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_5_rsc_req_obj_bcwt <= ~((~(din_5_rsc_req_obj_bcwt | din_5_rsc_req_obj_biwt))
          | din_5_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj_din_5_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj_din_5_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_5_rsc_req_obj_oswt, din_5_rsc_req_obj_vd, din_5_rsc_req_obj_biwt,
      din_5_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_5_rsc_req_obj_oswt;
  input din_5_rsc_req_obj_vd;
  output din_5_rsc_req_obj_biwt;
  output din_5_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_5_rsc_req_obj_pdswt0;
  reg din_5_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_5_rsc_req_obj_pdswt0 = (~ core_wten) & din_5_rsc_req_obj_oswt;
  assign din_5_rsc_req_obj_biwt = (din_5_rsc_req_obj_pdswt0 | din_5_rsc_req_obj_icwt)
      & din_5_rsc_req_obj_vd;
  assign din_5_rsc_req_obj_bdwt = din_5_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_5_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_5_rsc_req_obj_icwt <= ~((~(din_5_rsc_req_obj_icwt | din_5_rsc_req_obj_pdswt0))
          | din_5_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj_din_6_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj_din_6_rsc_req_wait_dp
    (
  clk, rst, din_6_rsc_req_obj_oswt, din_6_rsc_req_obj_wen_comp, din_6_rsc_req_obj_biwt,
      din_6_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_6_rsc_req_obj_oswt;
  output din_6_rsc_req_obj_wen_comp;
  input din_6_rsc_req_obj_biwt;
  input din_6_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_6_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_6_rsc_req_obj_wen_comp = (~ din_6_rsc_req_obj_oswt) | din_6_rsc_req_obj_biwt
      | din_6_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_6_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_6_rsc_req_obj_bcwt <= ~((~(din_6_rsc_req_obj_bcwt | din_6_rsc_req_obj_biwt))
          | din_6_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj_din_6_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj_din_6_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_6_rsc_req_obj_oswt, din_6_rsc_req_obj_vd, din_6_rsc_req_obj_biwt,
      din_6_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_6_rsc_req_obj_oswt;
  input din_6_rsc_req_obj_vd;
  output din_6_rsc_req_obj_biwt;
  output din_6_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_6_rsc_req_obj_pdswt0;
  reg din_6_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_6_rsc_req_obj_pdswt0 = (~ core_wten) & din_6_rsc_req_obj_oswt;
  assign din_6_rsc_req_obj_biwt = (din_6_rsc_req_obj_pdswt0 | din_6_rsc_req_obj_icwt)
      & din_6_rsc_req_obj_vd;
  assign din_6_rsc_req_obj_bdwt = din_6_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_6_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_6_rsc_req_obj_icwt <= ~((~(din_6_rsc_req_obj_icwt | din_6_rsc_req_obj_pdswt0))
          | din_6_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj_din_7_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj_din_7_rsc_req_wait_dp
    (
  clk, rst, din_7_rsc_req_obj_oswt, din_7_rsc_req_obj_wen_comp, din_7_rsc_req_obj_biwt,
      din_7_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_7_rsc_req_obj_oswt;
  output din_7_rsc_req_obj_wen_comp;
  input din_7_rsc_req_obj_biwt;
  input din_7_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_7_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_7_rsc_req_obj_wen_comp = (~ din_7_rsc_req_obj_oswt) | din_7_rsc_req_obj_biwt
      | din_7_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_7_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_7_rsc_req_obj_bcwt <= ~((~(din_7_rsc_req_obj_bcwt | din_7_rsc_req_obj_biwt))
          | din_7_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj_din_7_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj_din_7_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_7_rsc_req_obj_oswt, din_7_rsc_req_obj_vd, din_7_rsc_req_obj_biwt,
      din_7_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_7_rsc_req_obj_oswt;
  input din_7_rsc_req_obj_vd;
  output din_7_rsc_req_obj_biwt;
  output din_7_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_7_rsc_req_obj_pdswt0;
  reg din_7_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_7_rsc_req_obj_pdswt0 = (~ core_wten) & din_7_rsc_req_obj_oswt;
  assign din_7_rsc_req_obj_biwt = (din_7_rsc_req_obj_pdswt0 | din_7_rsc_req_obj_icwt)
      & din_7_rsc_req_obj_vd;
  assign din_7_rsc_req_obj_bdwt = din_7_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_7_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_7_rsc_req_obj_icwt <= ~((~(din_7_rsc_req_obj_icwt | din_7_rsc_req_obj_pdswt0))
          | din_7_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj_din_8_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj_din_8_rsc_req_wait_dp
    (
  clk, rst, din_8_rsc_req_obj_oswt, din_8_rsc_req_obj_wen_comp, din_8_rsc_req_obj_biwt,
      din_8_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_8_rsc_req_obj_oswt;
  output din_8_rsc_req_obj_wen_comp;
  input din_8_rsc_req_obj_biwt;
  input din_8_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_8_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_8_rsc_req_obj_wen_comp = (~ din_8_rsc_req_obj_oswt) | din_8_rsc_req_obj_biwt
      | din_8_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_8_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_8_rsc_req_obj_bcwt <= ~((~(din_8_rsc_req_obj_bcwt | din_8_rsc_req_obj_biwt))
          | din_8_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj_din_8_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj_din_8_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_8_rsc_req_obj_oswt, din_8_rsc_req_obj_vd, din_8_rsc_req_obj_biwt,
      din_8_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_8_rsc_req_obj_oswt;
  input din_8_rsc_req_obj_vd;
  output din_8_rsc_req_obj_biwt;
  output din_8_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_8_rsc_req_obj_pdswt0;
  reg din_8_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_8_rsc_req_obj_pdswt0 = (~ core_wten) & din_8_rsc_req_obj_oswt;
  assign din_8_rsc_req_obj_biwt = (din_8_rsc_req_obj_pdswt0 | din_8_rsc_req_obj_icwt)
      & din_8_rsc_req_obj_vd;
  assign din_8_rsc_req_obj_bdwt = din_8_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_8_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_8_rsc_req_obj_icwt <= ~((~(din_8_rsc_req_obj_icwt | din_8_rsc_req_obj_pdswt0))
          | din_8_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj_din_9_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj_din_9_rsc_req_wait_dp
    (
  clk, rst, din_9_rsc_req_obj_oswt, din_9_rsc_req_obj_wen_comp, din_9_rsc_req_obj_biwt,
      din_9_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_9_rsc_req_obj_oswt;
  output din_9_rsc_req_obj_wen_comp;
  input din_9_rsc_req_obj_biwt;
  input din_9_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_9_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_9_rsc_req_obj_wen_comp = (~ din_9_rsc_req_obj_oswt) | din_9_rsc_req_obj_biwt
      | din_9_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_9_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_9_rsc_req_obj_bcwt <= ~((~(din_9_rsc_req_obj_bcwt | din_9_rsc_req_obj_biwt))
          | din_9_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj_din_9_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj_din_9_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_9_rsc_req_obj_oswt, din_9_rsc_req_obj_vd, din_9_rsc_req_obj_biwt,
      din_9_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_9_rsc_req_obj_oswt;
  input din_9_rsc_req_obj_vd;
  output din_9_rsc_req_obj_biwt;
  output din_9_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_9_rsc_req_obj_pdswt0;
  reg din_9_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_9_rsc_req_obj_pdswt0 = (~ core_wten) & din_9_rsc_req_obj_oswt;
  assign din_9_rsc_req_obj_biwt = (din_9_rsc_req_obj_pdswt0 | din_9_rsc_req_obj_icwt)
      & din_9_rsc_req_obj_vd;
  assign din_9_rsc_req_obj_bdwt = din_9_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_9_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_9_rsc_req_obj_icwt <= ~((~(din_9_rsc_req_obj_icwt | din_9_rsc_req_obj_pdswt0))
          | din_9_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj_din_10_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj_din_10_rsc_req_wait_dp
    (
  clk, rst, din_10_rsc_req_obj_oswt, din_10_rsc_req_obj_wen_comp, din_10_rsc_req_obj_biwt,
      din_10_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_10_rsc_req_obj_oswt;
  output din_10_rsc_req_obj_wen_comp;
  input din_10_rsc_req_obj_biwt;
  input din_10_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_10_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_10_rsc_req_obj_wen_comp = (~ din_10_rsc_req_obj_oswt) | din_10_rsc_req_obj_biwt
      | din_10_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_10_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_10_rsc_req_obj_bcwt <= ~((~(din_10_rsc_req_obj_bcwt | din_10_rsc_req_obj_biwt))
          | din_10_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj_din_10_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj_din_10_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_10_rsc_req_obj_oswt, din_10_rsc_req_obj_vd,
      din_10_rsc_req_obj_biwt, din_10_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_10_rsc_req_obj_oswt;
  input din_10_rsc_req_obj_vd;
  output din_10_rsc_req_obj_biwt;
  output din_10_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_10_rsc_req_obj_pdswt0;
  reg din_10_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_10_rsc_req_obj_pdswt0 = (~ core_wten) & din_10_rsc_req_obj_oswt;
  assign din_10_rsc_req_obj_biwt = (din_10_rsc_req_obj_pdswt0 | din_10_rsc_req_obj_icwt)
      & din_10_rsc_req_obj_vd;
  assign din_10_rsc_req_obj_bdwt = din_10_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_10_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_10_rsc_req_obj_icwt <= ~((~(din_10_rsc_req_obj_icwt | din_10_rsc_req_obj_pdswt0))
          | din_10_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj_din_11_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj_din_11_rsc_req_wait_dp
    (
  clk, rst, din_11_rsc_req_obj_oswt, din_11_rsc_req_obj_wen_comp, din_11_rsc_req_obj_biwt,
      din_11_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_11_rsc_req_obj_oswt;
  output din_11_rsc_req_obj_wen_comp;
  input din_11_rsc_req_obj_biwt;
  input din_11_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_11_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_11_rsc_req_obj_wen_comp = (~ din_11_rsc_req_obj_oswt) | din_11_rsc_req_obj_biwt
      | din_11_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_11_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_11_rsc_req_obj_bcwt <= ~((~(din_11_rsc_req_obj_bcwt | din_11_rsc_req_obj_biwt))
          | din_11_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj_din_11_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj_din_11_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_11_rsc_req_obj_oswt, din_11_rsc_req_obj_vd,
      din_11_rsc_req_obj_biwt, din_11_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_11_rsc_req_obj_oswt;
  input din_11_rsc_req_obj_vd;
  output din_11_rsc_req_obj_biwt;
  output din_11_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_11_rsc_req_obj_pdswt0;
  reg din_11_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_11_rsc_req_obj_pdswt0 = (~ core_wten) & din_11_rsc_req_obj_oswt;
  assign din_11_rsc_req_obj_biwt = (din_11_rsc_req_obj_pdswt0 | din_11_rsc_req_obj_icwt)
      & din_11_rsc_req_obj_vd;
  assign din_11_rsc_req_obj_bdwt = din_11_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_11_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_11_rsc_req_obj_icwt <= ~((~(din_11_rsc_req_obj_icwt | din_11_rsc_req_obj_pdswt0))
          | din_11_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj_din_12_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj_din_12_rsc_req_wait_dp
    (
  clk, rst, din_12_rsc_req_obj_oswt, din_12_rsc_req_obj_wen_comp, din_12_rsc_req_obj_biwt,
      din_12_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_12_rsc_req_obj_oswt;
  output din_12_rsc_req_obj_wen_comp;
  input din_12_rsc_req_obj_biwt;
  input din_12_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_12_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_12_rsc_req_obj_wen_comp = (~ din_12_rsc_req_obj_oswt) | din_12_rsc_req_obj_biwt
      | din_12_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_12_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_12_rsc_req_obj_bcwt <= ~((~(din_12_rsc_req_obj_bcwt | din_12_rsc_req_obj_biwt))
          | din_12_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj_din_12_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj_din_12_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_12_rsc_req_obj_oswt, din_12_rsc_req_obj_vd,
      din_12_rsc_req_obj_biwt, din_12_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_12_rsc_req_obj_oswt;
  input din_12_rsc_req_obj_vd;
  output din_12_rsc_req_obj_biwt;
  output din_12_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_12_rsc_req_obj_pdswt0;
  reg din_12_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_12_rsc_req_obj_pdswt0 = (~ core_wten) & din_12_rsc_req_obj_oswt;
  assign din_12_rsc_req_obj_biwt = (din_12_rsc_req_obj_pdswt0 | din_12_rsc_req_obj_icwt)
      & din_12_rsc_req_obj_vd;
  assign din_12_rsc_req_obj_bdwt = din_12_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_12_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_12_rsc_req_obj_icwt <= ~((~(din_12_rsc_req_obj_icwt | din_12_rsc_req_obj_pdswt0))
          | din_12_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj_din_13_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj_din_13_rsc_req_wait_dp
    (
  clk, rst, din_13_rsc_req_obj_oswt, din_13_rsc_req_obj_wen_comp, din_13_rsc_req_obj_biwt,
      din_13_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_13_rsc_req_obj_oswt;
  output din_13_rsc_req_obj_wen_comp;
  input din_13_rsc_req_obj_biwt;
  input din_13_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_13_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_13_rsc_req_obj_wen_comp = (~ din_13_rsc_req_obj_oswt) | din_13_rsc_req_obj_biwt
      | din_13_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_13_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_13_rsc_req_obj_bcwt <= ~((~(din_13_rsc_req_obj_bcwt | din_13_rsc_req_obj_biwt))
          | din_13_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj_din_13_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj_din_13_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_13_rsc_req_obj_oswt, din_13_rsc_req_obj_vd,
      din_13_rsc_req_obj_biwt, din_13_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_13_rsc_req_obj_oswt;
  input din_13_rsc_req_obj_vd;
  output din_13_rsc_req_obj_biwt;
  output din_13_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_13_rsc_req_obj_pdswt0;
  reg din_13_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_13_rsc_req_obj_pdswt0 = (~ core_wten) & din_13_rsc_req_obj_oswt;
  assign din_13_rsc_req_obj_biwt = (din_13_rsc_req_obj_pdswt0 | din_13_rsc_req_obj_icwt)
      & din_13_rsc_req_obj_vd;
  assign din_13_rsc_req_obj_bdwt = din_13_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_13_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_13_rsc_req_obj_icwt <= ~((~(din_13_rsc_req_obj_icwt | din_13_rsc_req_obj_pdswt0))
          | din_13_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj_din_14_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj_din_14_rsc_req_wait_dp
    (
  clk, rst, din_14_rsc_req_obj_oswt, din_14_rsc_req_obj_wen_comp, din_14_rsc_req_obj_biwt,
      din_14_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_14_rsc_req_obj_oswt;
  output din_14_rsc_req_obj_wen_comp;
  input din_14_rsc_req_obj_biwt;
  input din_14_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_14_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_14_rsc_req_obj_wen_comp = (~ din_14_rsc_req_obj_oswt) | din_14_rsc_req_obj_biwt
      | din_14_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_14_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_14_rsc_req_obj_bcwt <= ~((~(din_14_rsc_req_obj_bcwt | din_14_rsc_req_obj_biwt))
          | din_14_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj_din_14_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj_din_14_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_14_rsc_req_obj_oswt, din_14_rsc_req_obj_vd,
      din_14_rsc_req_obj_biwt, din_14_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_14_rsc_req_obj_oswt;
  input din_14_rsc_req_obj_vd;
  output din_14_rsc_req_obj_biwt;
  output din_14_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_14_rsc_req_obj_pdswt0;
  reg din_14_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_14_rsc_req_obj_pdswt0 = (~ core_wten) & din_14_rsc_req_obj_oswt;
  assign din_14_rsc_req_obj_biwt = (din_14_rsc_req_obj_pdswt0 | din_14_rsc_req_obj_icwt)
      & din_14_rsc_req_obj_vd;
  assign din_14_rsc_req_obj_bdwt = din_14_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_14_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_14_rsc_req_obj_icwt <= ~((~(din_14_rsc_req_obj_icwt | din_14_rsc_req_obj_pdswt0))
          | din_14_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj_din_15_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj_din_15_rsc_req_wait_dp
    (
  clk, rst, din_15_rsc_req_obj_oswt, din_15_rsc_req_obj_wen_comp, din_15_rsc_req_obj_biwt,
      din_15_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_15_rsc_req_obj_oswt;
  output din_15_rsc_req_obj_wen_comp;
  input din_15_rsc_req_obj_biwt;
  input din_15_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_15_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_15_rsc_req_obj_wen_comp = (~ din_15_rsc_req_obj_oswt) | din_15_rsc_req_obj_biwt
      | din_15_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_15_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_15_rsc_req_obj_bcwt <= ~((~(din_15_rsc_req_obj_bcwt | din_15_rsc_req_obj_biwt))
          | din_15_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj_din_15_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj_din_15_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_15_rsc_req_obj_oswt, din_15_rsc_req_obj_vd,
      din_15_rsc_req_obj_biwt, din_15_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_15_rsc_req_obj_oswt;
  input din_15_rsc_req_obj_vd;
  output din_15_rsc_req_obj_biwt;
  output din_15_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_15_rsc_req_obj_pdswt0;
  reg din_15_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_15_rsc_req_obj_pdswt0 = (~ core_wten) & din_15_rsc_req_obj_oswt;
  assign din_15_rsc_req_obj_biwt = (din_15_rsc_req_obj_pdswt0 | din_15_rsc_req_obj_icwt)
      & din_15_rsc_req_obj_vd;
  assign din_15_rsc_req_obj_bdwt = din_15_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_15_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_15_rsc_req_obj_icwt <= ~((~(din_15_rsc_req_obj_icwt | din_15_rsc_req_obj_pdswt0))
          | din_15_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj_din_16_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj_din_16_rsc_req_wait_dp
    (
  clk, rst, din_16_rsc_req_obj_oswt, din_16_rsc_req_obj_wen_comp, din_16_rsc_req_obj_biwt,
      din_16_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_16_rsc_req_obj_oswt;
  output din_16_rsc_req_obj_wen_comp;
  input din_16_rsc_req_obj_biwt;
  input din_16_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_16_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_16_rsc_req_obj_wen_comp = (~ din_16_rsc_req_obj_oswt) | din_16_rsc_req_obj_biwt
      | din_16_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_16_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_16_rsc_req_obj_bcwt <= ~((~(din_16_rsc_req_obj_bcwt | din_16_rsc_req_obj_biwt))
          | din_16_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj_din_16_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj_din_16_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_16_rsc_req_obj_oswt, din_16_rsc_req_obj_vd,
      din_16_rsc_req_obj_biwt, din_16_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_16_rsc_req_obj_oswt;
  input din_16_rsc_req_obj_vd;
  output din_16_rsc_req_obj_biwt;
  output din_16_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_16_rsc_req_obj_pdswt0;
  reg din_16_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_16_rsc_req_obj_pdswt0 = (~ core_wten) & din_16_rsc_req_obj_oswt;
  assign din_16_rsc_req_obj_biwt = (din_16_rsc_req_obj_pdswt0 | din_16_rsc_req_obj_icwt)
      & din_16_rsc_req_obj_vd;
  assign din_16_rsc_req_obj_bdwt = din_16_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_16_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_16_rsc_req_obj_icwt <= ~((~(din_16_rsc_req_obj_icwt | din_16_rsc_req_obj_pdswt0))
          | din_16_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj_din_17_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj_din_17_rsc_req_wait_dp
    (
  clk, rst, din_17_rsc_req_obj_oswt, din_17_rsc_req_obj_wen_comp, din_17_rsc_req_obj_biwt,
      din_17_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_17_rsc_req_obj_oswt;
  output din_17_rsc_req_obj_wen_comp;
  input din_17_rsc_req_obj_biwt;
  input din_17_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_17_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_17_rsc_req_obj_wen_comp = (~ din_17_rsc_req_obj_oswt) | din_17_rsc_req_obj_biwt
      | din_17_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_17_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_17_rsc_req_obj_bcwt <= ~((~(din_17_rsc_req_obj_bcwt | din_17_rsc_req_obj_biwt))
          | din_17_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj_din_17_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj_din_17_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_17_rsc_req_obj_oswt, din_17_rsc_req_obj_vd,
      din_17_rsc_req_obj_biwt, din_17_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_17_rsc_req_obj_oswt;
  input din_17_rsc_req_obj_vd;
  output din_17_rsc_req_obj_biwt;
  output din_17_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_17_rsc_req_obj_pdswt0;
  reg din_17_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_17_rsc_req_obj_pdswt0 = (~ core_wten) & din_17_rsc_req_obj_oswt;
  assign din_17_rsc_req_obj_biwt = (din_17_rsc_req_obj_pdswt0 | din_17_rsc_req_obj_icwt)
      & din_17_rsc_req_obj_vd;
  assign din_17_rsc_req_obj_bdwt = din_17_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_17_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_17_rsc_req_obj_icwt <= ~((~(din_17_rsc_req_obj_icwt | din_17_rsc_req_obj_pdswt0))
          | din_17_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_rls_obj_din_17_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_rls_obj_din_17_rsc_rls_wait_ctrl
    (
  core_wten, din_17_rsc_rls_obj_iswt0, din_17_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_17_rsc_rls_obj_iswt0;
  output din_17_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_17_rsc_rls_obj_ld_core_sct = din_17_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_rls_obj_din_16_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_rls_obj_din_16_rsc_rls_wait_ctrl
    (
  core_wten, din_16_rsc_rls_obj_iswt0, din_16_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_16_rsc_rls_obj_iswt0;
  output din_16_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_16_rsc_rls_obj_ld_core_sct = din_16_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_rls_obj_din_15_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_rls_obj_din_15_rsc_rls_wait_ctrl
    (
  core_wten, din_15_rsc_rls_obj_iswt0, din_15_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_15_rsc_rls_obj_iswt0;
  output din_15_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_15_rsc_rls_obj_ld_core_sct = din_15_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_rls_obj_din_14_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_rls_obj_din_14_rsc_rls_wait_ctrl
    (
  core_wten, din_14_rsc_rls_obj_iswt0, din_14_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_14_rsc_rls_obj_iswt0;
  output din_14_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_14_rsc_rls_obj_ld_core_sct = din_14_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_rls_obj_din_13_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_rls_obj_din_13_rsc_rls_wait_ctrl
    (
  core_wten, din_13_rsc_rls_obj_iswt0, din_13_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_13_rsc_rls_obj_iswt0;
  output din_13_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_13_rsc_rls_obj_ld_core_sct = din_13_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_rls_obj_din_12_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_rls_obj_din_12_rsc_rls_wait_ctrl
    (
  core_wten, din_12_rsc_rls_obj_iswt0, din_12_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_12_rsc_rls_obj_iswt0;
  output din_12_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_12_rsc_rls_obj_ld_core_sct = din_12_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_rls_obj_din_11_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_rls_obj_din_11_rsc_rls_wait_ctrl
    (
  core_wten, din_11_rsc_rls_obj_iswt0, din_11_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_11_rsc_rls_obj_iswt0;
  output din_11_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_11_rsc_rls_obj_ld_core_sct = din_11_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_rls_obj_din_10_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_rls_obj_din_10_rsc_rls_wait_ctrl
    (
  core_wten, din_10_rsc_rls_obj_iswt0, din_10_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_10_rsc_rls_obj_iswt0;
  output din_10_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_10_rsc_rls_obj_ld_core_sct = din_10_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_rls_obj_din_9_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_rls_obj_din_9_rsc_rls_wait_ctrl
    (
  core_wten, din_9_rsc_rls_obj_iswt0, din_9_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_9_rsc_rls_obj_iswt0;
  output din_9_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_9_rsc_rls_obj_ld_core_sct = din_9_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_rls_obj_din_8_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_rls_obj_din_8_rsc_rls_wait_ctrl
    (
  core_wten, din_8_rsc_rls_obj_iswt0, din_8_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_8_rsc_rls_obj_iswt0;
  output din_8_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_8_rsc_rls_obj_ld_core_sct = din_8_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_rls_obj_din_7_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_rls_obj_din_7_rsc_rls_wait_ctrl
    (
  core_wten, din_7_rsc_rls_obj_iswt0, din_7_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_7_rsc_rls_obj_iswt0;
  output din_7_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_7_rsc_rls_obj_ld_core_sct = din_7_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_rls_obj_din_6_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_rls_obj_din_6_rsc_rls_wait_ctrl
    (
  core_wten, din_6_rsc_rls_obj_iswt0, din_6_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_6_rsc_rls_obj_iswt0;
  output din_6_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_6_rsc_rls_obj_ld_core_sct = din_6_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_rls_obj_din_5_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_rls_obj_din_5_rsc_rls_wait_ctrl
    (
  core_wten, din_5_rsc_rls_obj_iswt0, din_5_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_5_rsc_rls_obj_iswt0;
  output din_5_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_5_rsc_rls_obj_ld_core_sct = din_5_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_rls_obj_din_4_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_rls_obj_din_4_rsc_rls_wait_ctrl
    (
  core_wten, din_4_rsc_rls_obj_iswt0, din_4_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_4_rsc_rls_obj_iswt0;
  output din_4_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_4_rsc_rls_obj_ld_core_sct = din_4_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_rls_obj_din_3_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_rls_obj_din_3_rsc_rls_wait_ctrl
    (
  core_wten, din_3_rsc_rls_obj_iswt0, din_3_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_3_rsc_rls_obj_iswt0;
  output din_3_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_3_rsc_rls_obj_ld_core_sct = din_3_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_rls_obj_din_2_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_rls_obj_din_2_rsc_rls_wait_ctrl
    (
  core_wten, din_2_rsc_rls_obj_iswt0, din_2_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_2_rsc_rls_obj_iswt0;
  output din_2_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_2_rsc_rls_obj_ld_core_sct = din_2_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_rls_obj_din_1_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_rls_obj_din_1_rsc_rls_wait_ctrl
    (
  core_wten, din_1_rsc_rls_obj_iswt0, din_1_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_1_rsc_rls_obj_iswt0;
  output din_1_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_1_rsc_rls_obj_ld_core_sct = din_1_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_rls_obj_din_0_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_rls_obj_din_0_rsc_rls_wait_ctrl
    (
  core_wten, din_0_rsc_rls_obj_iswt0, din_0_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_0_rsc_rls_obj_iswt0;
  output din_0_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_0_rsc_rls_obj_ld_core_sct = din_0_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_dout_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_dout_wait_dp (
  clk, rst, dout_rsci_oswt, dout_rsci_wen_comp, dout_rsci_biwt, dout_rsci_bdwt
);
  input clk;
  input rst;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input dout_rsci_biwt;
  input dout_rsci_bdwt;


  // Interconnect Declarations
  reg dout_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_wen_comp = (~ dout_rsci_oswt) | dout_rsci_biwt | dout_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_bcwt <= 1'b0;
    end
    else begin
      dout_rsci_bcwt <= ~((~(dout_rsci_bcwt | dout_rsci_biwt)) | dout_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_dout_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_dout_wait_ctrl (
  clk, rst, core_wen, core_wten, dout_rsci_oswt, dout_rsci_biwt, dout_rsci_bdwt,
      dout_rsci_ld_core_sct, dout_rsci_vd
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_rsci_oswt;
  output dout_rsci_biwt;
  output dout_rsci_bdwt;
  output dout_rsci_ld_core_sct;
  input dout_rsci_vd;


  // Interconnect Declarations
  wire dout_rsci_ogwt;
  wire dout_rsci_pdswt0;
  reg dout_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_pdswt0 = (~ core_wten) & dout_rsci_oswt;
  assign dout_rsci_biwt = dout_rsci_ogwt & dout_rsci_vd;
  assign dout_rsci_ogwt = dout_rsci_pdswt0 | dout_rsci_icwt;
  assign dout_rsci_bdwt = dout_rsci_oswt & core_wen;
  assign dout_rsci_ld_core_sct = dout_rsci_oswt & dout_rsci_ogwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_icwt <= 1'b0;
    end
    else begin
      dout_rsci_icwt <= ~((~(dout_rsci_icwt | dout_rsci_pdswt0)) | dout_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1_din_17_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1_din_17_rsc_wait_dp (
  clk, rst, din_17_rsci_douta_d, din_17_rsci_douta_d_mxwt, din_17_rsci_biwt, din_17_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_17_rsci_douta_d;
  output [15:0] din_17_rsci_douta_d_mxwt;
  input din_17_rsci_biwt;
  input din_17_rsci_bdwt;


  // Interconnect Declarations
  reg din_17_rsci_bcwt;
  reg [15:0] din_17_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_17_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_17_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_17_rsci_douta_d[15:0]),
      din_17_rsci_douta_d_bfwt_15_0, din_17_rsci_bcwt);
  assign din_17_rsci_douta_d_mxwt = din_17_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_17_rsci_bcwt <= 1'b0;
      din_17_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_17_rsci_bcwt <= ~((~(din_17_rsci_bcwt | din_17_rsci_biwt)) | din_17_rsci_bdwt);
      din_17_rsci_douta_d_bfwt_15_0 <= din_17_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1_din_17_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1_din_17_rsc_wait_ctrl
    (
  core_wen, core_wten, din_17_rsci_oswt, din_17_rsci_biwt, din_17_rsci_bdwt, din_17_rsci_biwt_pff,
      din_17_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_17_rsci_oswt;
  output din_17_rsci_biwt;
  output din_17_rsci_bdwt;
  output din_17_rsci_biwt_pff;
  input din_17_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_17_rsci_bdwt = din_17_rsci_oswt & core_wen;
  assign din_17_rsci_biwt = (~ core_wten) & din_17_rsci_oswt;
  assign din_17_rsci_biwt_pff = core_wen & din_17_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1_din_16_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1_din_16_rsc_wait_dp (
  clk, rst, din_16_rsci_douta_d, din_16_rsci_douta_d_mxwt, din_16_rsci_biwt, din_16_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_16_rsci_douta_d;
  output [15:0] din_16_rsci_douta_d_mxwt;
  input din_16_rsci_biwt;
  input din_16_rsci_bdwt;


  // Interconnect Declarations
  reg din_16_rsci_bcwt;
  reg [15:0] din_16_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_16_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_16_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_16_rsci_douta_d[15:0]),
      din_16_rsci_douta_d_bfwt_15_0, din_16_rsci_bcwt);
  assign din_16_rsci_douta_d_mxwt = din_16_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_16_rsci_bcwt <= 1'b0;
      din_16_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_16_rsci_bcwt <= ~((~(din_16_rsci_bcwt | din_16_rsci_biwt)) | din_16_rsci_bdwt);
      din_16_rsci_douta_d_bfwt_15_0 <= din_16_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1_din_16_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1_din_16_rsc_wait_ctrl
    (
  core_wen, core_wten, din_16_rsci_oswt, din_16_rsci_biwt, din_16_rsci_bdwt, din_16_rsci_biwt_pff,
      din_16_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_16_rsci_oswt;
  output din_16_rsci_biwt;
  output din_16_rsci_bdwt;
  output din_16_rsci_biwt_pff;
  input din_16_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_16_rsci_bdwt = din_16_rsci_oswt & core_wen;
  assign din_16_rsci_biwt = (~ core_wten) & din_16_rsci_oswt;
  assign din_16_rsci_biwt_pff = core_wen & din_16_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1_din_15_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1_din_15_rsc_wait_dp (
  clk, rst, din_15_rsci_douta_d, din_15_rsci_douta_d_mxwt, din_15_rsci_biwt, din_15_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_15_rsci_douta_d;
  output [15:0] din_15_rsci_douta_d_mxwt;
  input din_15_rsci_biwt;
  input din_15_rsci_bdwt;


  // Interconnect Declarations
  reg din_15_rsci_bcwt;
  reg [15:0] din_15_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_15_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_15_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_15_rsci_douta_d[15:0]),
      din_15_rsci_douta_d_bfwt_15_0, din_15_rsci_bcwt);
  assign din_15_rsci_douta_d_mxwt = din_15_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_15_rsci_bcwt <= 1'b0;
      din_15_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_15_rsci_bcwt <= ~((~(din_15_rsci_bcwt | din_15_rsci_biwt)) | din_15_rsci_bdwt);
      din_15_rsci_douta_d_bfwt_15_0 <= din_15_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1_din_15_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1_din_15_rsc_wait_ctrl
    (
  core_wen, core_wten, din_15_rsci_oswt, din_15_rsci_biwt, din_15_rsci_bdwt, din_15_rsci_biwt_pff,
      din_15_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_15_rsci_oswt;
  output din_15_rsci_biwt;
  output din_15_rsci_bdwt;
  output din_15_rsci_biwt_pff;
  input din_15_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_15_rsci_bdwt = din_15_rsci_oswt & core_wen;
  assign din_15_rsci_biwt = (~ core_wten) & din_15_rsci_oswt;
  assign din_15_rsci_biwt_pff = core_wen & din_15_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1_din_14_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1_din_14_rsc_wait_dp (
  clk, rst, din_14_rsci_douta_d, din_14_rsci_douta_d_mxwt, din_14_rsci_biwt, din_14_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_14_rsci_douta_d;
  output [15:0] din_14_rsci_douta_d_mxwt;
  input din_14_rsci_biwt;
  input din_14_rsci_bdwt;


  // Interconnect Declarations
  reg din_14_rsci_bcwt;
  reg [15:0] din_14_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_14_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_14_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_14_rsci_douta_d[15:0]),
      din_14_rsci_douta_d_bfwt_15_0, din_14_rsci_bcwt);
  assign din_14_rsci_douta_d_mxwt = din_14_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_14_rsci_bcwt <= 1'b0;
      din_14_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_14_rsci_bcwt <= ~((~(din_14_rsci_bcwt | din_14_rsci_biwt)) | din_14_rsci_bdwt);
      din_14_rsci_douta_d_bfwt_15_0 <= din_14_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1_din_14_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1_din_14_rsc_wait_ctrl
    (
  core_wen, core_wten, din_14_rsci_oswt, din_14_rsci_biwt, din_14_rsci_bdwt, din_14_rsci_biwt_pff,
      din_14_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_14_rsci_oswt;
  output din_14_rsci_biwt;
  output din_14_rsci_bdwt;
  output din_14_rsci_biwt_pff;
  input din_14_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_14_rsci_bdwt = din_14_rsci_oswt & core_wen;
  assign din_14_rsci_biwt = (~ core_wten) & din_14_rsci_oswt;
  assign din_14_rsci_biwt_pff = core_wen & din_14_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1_din_13_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1_din_13_rsc_wait_dp (
  clk, rst, din_13_rsci_douta_d, din_13_rsci_douta_d_mxwt, din_13_rsci_biwt, din_13_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_13_rsci_douta_d;
  output [15:0] din_13_rsci_douta_d_mxwt;
  input din_13_rsci_biwt;
  input din_13_rsci_bdwt;


  // Interconnect Declarations
  reg din_13_rsci_bcwt;
  reg [15:0] din_13_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_13_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_13_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_13_rsci_douta_d[15:0]),
      din_13_rsci_douta_d_bfwt_15_0, din_13_rsci_bcwt);
  assign din_13_rsci_douta_d_mxwt = din_13_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_13_rsci_bcwt <= 1'b0;
      din_13_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_13_rsci_bcwt <= ~((~(din_13_rsci_bcwt | din_13_rsci_biwt)) | din_13_rsci_bdwt);
      din_13_rsci_douta_d_bfwt_15_0 <= din_13_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1_din_13_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1_din_13_rsc_wait_ctrl
    (
  core_wen, core_wten, din_13_rsci_oswt, din_13_rsci_biwt, din_13_rsci_bdwt, din_13_rsci_biwt_pff,
      din_13_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_13_rsci_oswt;
  output din_13_rsci_biwt;
  output din_13_rsci_bdwt;
  output din_13_rsci_biwt_pff;
  input din_13_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_13_rsci_bdwt = din_13_rsci_oswt & core_wen;
  assign din_13_rsci_biwt = (~ core_wten) & din_13_rsci_oswt;
  assign din_13_rsci_biwt_pff = core_wen & din_13_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1_din_12_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1_din_12_rsc_wait_dp (
  clk, rst, din_12_rsci_douta_d, din_12_rsci_douta_d_mxwt, din_12_rsci_biwt, din_12_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_12_rsci_douta_d;
  output [15:0] din_12_rsci_douta_d_mxwt;
  input din_12_rsci_biwt;
  input din_12_rsci_bdwt;


  // Interconnect Declarations
  reg din_12_rsci_bcwt;
  reg [15:0] din_12_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_12_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_12_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_12_rsci_douta_d[15:0]),
      din_12_rsci_douta_d_bfwt_15_0, din_12_rsci_bcwt);
  assign din_12_rsci_douta_d_mxwt = din_12_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_12_rsci_bcwt <= 1'b0;
      din_12_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_12_rsci_bcwt <= ~((~(din_12_rsci_bcwt | din_12_rsci_biwt)) | din_12_rsci_bdwt);
      din_12_rsci_douta_d_bfwt_15_0 <= din_12_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1_din_12_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1_din_12_rsc_wait_ctrl
    (
  core_wen, core_wten, din_12_rsci_oswt, din_12_rsci_biwt, din_12_rsci_bdwt, din_12_rsci_biwt_pff,
      din_12_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_12_rsci_oswt;
  output din_12_rsci_biwt;
  output din_12_rsci_bdwt;
  output din_12_rsci_biwt_pff;
  input din_12_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_12_rsci_bdwt = din_12_rsci_oswt & core_wen;
  assign din_12_rsci_biwt = (~ core_wten) & din_12_rsci_oswt;
  assign din_12_rsci_biwt_pff = core_wen & din_12_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1_din_11_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1_din_11_rsc_wait_dp (
  clk, rst, din_11_rsci_douta_d, din_11_rsci_douta_d_mxwt, din_11_rsci_biwt, din_11_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_11_rsci_douta_d;
  output [15:0] din_11_rsci_douta_d_mxwt;
  input din_11_rsci_biwt;
  input din_11_rsci_bdwt;


  // Interconnect Declarations
  reg din_11_rsci_bcwt;
  reg [15:0] din_11_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_11_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_11_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_11_rsci_douta_d[15:0]),
      din_11_rsci_douta_d_bfwt_15_0, din_11_rsci_bcwt);
  assign din_11_rsci_douta_d_mxwt = din_11_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_11_rsci_bcwt <= 1'b0;
      din_11_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_11_rsci_bcwt <= ~((~(din_11_rsci_bcwt | din_11_rsci_biwt)) | din_11_rsci_bdwt);
      din_11_rsci_douta_d_bfwt_15_0 <= din_11_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1_din_11_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1_din_11_rsc_wait_ctrl
    (
  core_wen, core_wten, din_11_rsci_oswt, din_11_rsci_biwt, din_11_rsci_bdwt, din_11_rsci_biwt_pff,
      din_11_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_11_rsci_oswt;
  output din_11_rsci_biwt;
  output din_11_rsci_bdwt;
  output din_11_rsci_biwt_pff;
  input din_11_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_11_rsci_bdwt = din_11_rsci_oswt & core_wen;
  assign din_11_rsci_biwt = (~ core_wten) & din_11_rsci_oswt;
  assign din_11_rsci_biwt_pff = core_wen & din_11_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1_din_10_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1_din_10_rsc_wait_dp (
  clk, rst, din_10_rsci_douta_d, din_10_rsci_douta_d_mxwt, din_10_rsci_biwt, din_10_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_10_rsci_douta_d;
  output [15:0] din_10_rsci_douta_d_mxwt;
  input din_10_rsci_biwt;
  input din_10_rsci_bdwt;


  // Interconnect Declarations
  reg din_10_rsci_bcwt;
  reg [15:0] din_10_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_10_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_10_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_10_rsci_douta_d[15:0]),
      din_10_rsci_douta_d_bfwt_15_0, din_10_rsci_bcwt);
  assign din_10_rsci_douta_d_mxwt = din_10_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_10_rsci_bcwt <= 1'b0;
      din_10_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_10_rsci_bcwt <= ~((~(din_10_rsci_bcwt | din_10_rsci_biwt)) | din_10_rsci_bdwt);
      din_10_rsci_douta_d_bfwt_15_0 <= din_10_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1_din_10_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1_din_10_rsc_wait_ctrl
    (
  core_wen, core_wten, din_10_rsci_oswt, din_10_rsci_biwt, din_10_rsci_bdwt, din_10_rsci_biwt_pff,
      din_10_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_10_rsci_oswt;
  output din_10_rsci_biwt;
  output din_10_rsci_bdwt;
  output din_10_rsci_biwt_pff;
  input din_10_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_10_rsci_bdwt = din_10_rsci_oswt & core_wen;
  assign din_10_rsci_biwt = (~ core_wten) & din_10_rsci_oswt;
  assign din_10_rsci_biwt_pff = core_wen & din_10_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1_din_9_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1_din_9_rsc_wait_dp (
  clk, rst, din_9_rsci_douta_d, din_9_rsci_douta_d_mxwt, din_9_rsci_biwt, din_9_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_9_rsci_douta_d;
  output [15:0] din_9_rsci_douta_d_mxwt;
  input din_9_rsci_biwt;
  input din_9_rsci_bdwt;


  // Interconnect Declarations
  reg din_9_rsci_bcwt;
  reg [15:0] din_9_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_9_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_9_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_9_rsci_douta_d[15:0]),
      din_9_rsci_douta_d_bfwt_15_0, din_9_rsci_bcwt);
  assign din_9_rsci_douta_d_mxwt = din_9_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_9_rsci_bcwt <= 1'b0;
      din_9_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_9_rsci_bcwt <= ~((~(din_9_rsci_bcwt | din_9_rsci_biwt)) | din_9_rsci_bdwt);
      din_9_rsci_douta_d_bfwt_15_0 <= din_9_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1_din_9_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1_din_9_rsc_wait_ctrl (
  core_wen, core_wten, din_9_rsci_oswt, din_9_rsci_biwt, din_9_rsci_bdwt, din_9_rsci_biwt_pff,
      din_9_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_9_rsci_oswt;
  output din_9_rsci_biwt;
  output din_9_rsci_bdwt;
  output din_9_rsci_biwt_pff;
  input din_9_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_9_rsci_bdwt = din_9_rsci_oswt & core_wen;
  assign din_9_rsci_biwt = (~ core_wten) & din_9_rsci_oswt;
  assign din_9_rsci_biwt_pff = core_wen & din_9_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1_din_8_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1_din_8_rsc_wait_dp (
  clk, rst, din_8_rsci_douta_d, din_8_rsci_douta_d_mxwt, din_8_rsci_biwt, din_8_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_8_rsci_douta_d;
  output [15:0] din_8_rsci_douta_d_mxwt;
  input din_8_rsci_biwt;
  input din_8_rsci_bdwt;


  // Interconnect Declarations
  reg din_8_rsci_bcwt;
  reg [15:0] din_8_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_8_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_8_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_8_rsci_douta_d[15:0]),
      din_8_rsci_douta_d_bfwt_15_0, din_8_rsci_bcwt);
  assign din_8_rsci_douta_d_mxwt = din_8_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_8_rsci_bcwt <= 1'b0;
      din_8_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_8_rsci_bcwt <= ~((~(din_8_rsci_bcwt | din_8_rsci_biwt)) | din_8_rsci_bdwt);
      din_8_rsci_douta_d_bfwt_15_0 <= din_8_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1_din_8_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1_din_8_rsc_wait_ctrl (
  core_wen, core_wten, din_8_rsci_oswt, din_8_rsci_biwt, din_8_rsci_bdwt, din_8_rsci_biwt_pff,
      din_8_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_8_rsci_oswt;
  output din_8_rsci_biwt;
  output din_8_rsci_bdwt;
  output din_8_rsci_biwt_pff;
  input din_8_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_8_rsci_bdwt = din_8_rsci_oswt & core_wen;
  assign din_8_rsci_biwt = (~ core_wten) & din_8_rsci_oswt;
  assign din_8_rsci_biwt_pff = core_wen & din_8_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1_din_7_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1_din_7_rsc_wait_dp (
  clk, rst, din_7_rsci_douta_d, din_7_rsci_douta_d_mxwt, din_7_rsci_biwt, din_7_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_7_rsci_douta_d;
  output [15:0] din_7_rsci_douta_d_mxwt;
  input din_7_rsci_biwt;
  input din_7_rsci_bdwt;


  // Interconnect Declarations
  reg din_7_rsci_bcwt;
  reg [15:0] din_7_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_7_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_7_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_7_rsci_douta_d[15:0]),
      din_7_rsci_douta_d_bfwt_15_0, din_7_rsci_bcwt);
  assign din_7_rsci_douta_d_mxwt = din_7_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_7_rsci_bcwt <= 1'b0;
      din_7_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_7_rsci_bcwt <= ~((~(din_7_rsci_bcwt | din_7_rsci_biwt)) | din_7_rsci_bdwt);
      din_7_rsci_douta_d_bfwt_15_0 <= din_7_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1_din_7_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1_din_7_rsc_wait_ctrl (
  core_wen, core_wten, din_7_rsci_oswt, din_7_rsci_biwt, din_7_rsci_bdwt, din_7_rsci_biwt_pff,
      din_7_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_7_rsci_oswt;
  output din_7_rsci_biwt;
  output din_7_rsci_bdwt;
  output din_7_rsci_biwt_pff;
  input din_7_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_7_rsci_bdwt = din_7_rsci_oswt & core_wen;
  assign din_7_rsci_biwt = (~ core_wten) & din_7_rsci_oswt;
  assign din_7_rsci_biwt_pff = core_wen & din_7_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1_din_6_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1_din_6_rsc_wait_dp (
  clk, rst, din_6_rsci_douta_d, din_6_rsci_douta_d_mxwt, din_6_rsci_biwt, din_6_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_6_rsci_douta_d;
  output [15:0] din_6_rsci_douta_d_mxwt;
  input din_6_rsci_biwt;
  input din_6_rsci_bdwt;


  // Interconnect Declarations
  reg din_6_rsci_bcwt;
  reg [15:0] din_6_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_6_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_6_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_6_rsci_douta_d[15:0]),
      din_6_rsci_douta_d_bfwt_15_0, din_6_rsci_bcwt);
  assign din_6_rsci_douta_d_mxwt = din_6_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_6_rsci_bcwt <= 1'b0;
      din_6_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_6_rsci_bcwt <= ~((~(din_6_rsci_bcwt | din_6_rsci_biwt)) | din_6_rsci_bdwt);
      din_6_rsci_douta_d_bfwt_15_0 <= din_6_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1_din_6_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1_din_6_rsc_wait_ctrl (
  core_wen, core_wten, din_6_rsci_oswt, din_6_rsci_biwt, din_6_rsci_bdwt, din_6_rsci_biwt_pff,
      din_6_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_6_rsci_oswt;
  output din_6_rsci_biwt;
  output din_6_rsci_bdwt;
  output din_6_rsci_biwt_pff;
  input din_6_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_6_rsci_bdwt = din_6_rsci_oswt & core_wen;
  assign din_6_rsci_biwt = (~ core_wten) & din_6_rsci_oswt;
  assign din_6_rsci_biwt_pff = core_wen & din_6_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1_din_5_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1_din_5_rsc_wait_dp (
  clk, rst, din_5_rsci_douta_d, din_5_rsci_douta_d_mxwt, din_5_rsci_biwt, din_5_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_5_rsci_douta_d;
  output [15:0] din_5_rsci_douta_d_mxwt;
  input din_5_rsci_biwt;
  input din_5_rsci_bdwt;


  // Interconnect Declarations
  reg din_5_rsci_bcwt;
  reg [15:0] din_5_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_5_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_5_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_5_rsci_douta_d[15:0]),
      din_5_rsci_douta_d_bfwt_15_0, din_5_rsci_bcwt);
  assign din_5_rsci_douta_d_mxwt = din_5_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_5_rsci_bcwt <= 1'b0;
      din_5_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_5_rsci_bcwt <= ~((~(din_5_rsci_bcwt | din_5_rsci_biwt)) | din_5_rsci_bdwt);
      din_5_rsci_douta_d_bfwt_15_0 <= din_5_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1_din_5_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1_din_5_rsc_wait_ctrl (
  core_wen, core_wten, din_5_rsci_oswt, din_5_rsci_biwt, din_5_rsci_bdwt, din_5_rsci_biwt_pff,
      din_5_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_5_rsci_oswt;
  output din_5_rsci_biwt;
  output din_5_rsci_bdwt;
  output din_5_rsci_biwt_pff;
  input din_5_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_5_rsci_bdwt = din_5_rsci_oswt & core_wen;
  assign din_5_rsci_biwt = (~ core_wten) & din_5_rsci_oswt;
  assign din_5_rsci_biwt_pff = core_wen & din_5_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1_din_4_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1_din_4_rsc_wait_dp (
  clk, rst, din_4_rsci_douta_d, din_4_rsci_douta_d_mxwt, din_4_rsci_biwt, din_4_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_4_rsci_douta_d;
  output [15:0] din_4_rsci_douta_d_mxwt;
  input din_4_rsci_biwt;
  input din_4_rsci_bdwt;


  // Interconnect Declarations
  reg din_4_rsci_bcwt;
  reg [15:0] din_4_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_4_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_4_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_4_rsci_douta_d[15:0]),
      din_4_rsci_douta_d_bfwt_15_0, din_4_rsci_bcwt);
  assign din_4_rsci_douta_d_mxwt = din_4_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_4_rsci_bcwt <= 1'b0;
      din_4_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_4_rsci_bcwt <= ~((~(din_4_rsci_bcwt | din_4_rsci_biwt)) | din_4_rsci_bdwt);
      din_4_rsci_douta_d_bfwt_15_0 <= din_4_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1_din_4_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1_din_4_rsc_wait_ctrl (
  core_wen, core_wten, din_4_rsci_oswt, din_4_rsci_biwt, din_4_rsci_bdwt, din_4_rsci_biwt_pff,
      din_4_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_4_rsci_oswt;
  output din_4_rsci_biwt;
  output din_4_rsci_bdwt;
  output din_4_rsci_biwt_pff;
  input din_4_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_4_rsci_bdwt = din_4_rsci_oswt & core_wen;
  assign din_4_rsci_biwt = (~ core_wten) & din_4_rsci_oswt;
  assign din_4_rsci_biwt_pff = core_wen & din_4_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1_din_3_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1_din_3_rsc_wait_dp (
  clk, rst, din_3_rsci_douta_d, din_3_rsci_douta_d_mxwt, din_3_rsci_biwt, din_3_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_3_rsci_douta_d;
  output [15:0] din_3_rsci_douta_d_mxwt;
  input din_3_rsci_biwt;
  input din_3_rsci_bdwt;


  // Interconnect Declarations
  reg din_3_rsci_bcwt;
  reg [15:0] din_3_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_3_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_3_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_3_rsci_douta_d[15:0]),
      din_3_rsci_douta_d_bfwt_15_0, din_3_rsci_bcwt);
  assign din_3_rsci_douta_d_mxwt = din_3_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_3_rsci_bcwt <= 1'b0;
      din_3_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_3_rsci_bcwt <= ~((~(din_3_rsci_bcwt | din_3_rsci_biwt)) | din_3_rsci_bdwt);
      din_3_rsci_douta_d_bfwt_15_0 <= din_3_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1_din_3_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1_din_3_rsc_wait_ctrl (
  core_wen, core_wten, din_3_rsci_oswt, din_3_rsci_biwt, din_3_rsci_bdwt, din_3_rsci_biwt_pff,
      din_3_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_3_rsci_oswt;
  output din_3_rsci_biwt;
  output din_3_rsci_bdwt;
  output din_3_rsci_biwt_pff;
  input din_3_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_3_rsci_bdwt = din_3_rsci_oswt & core_wen;
  assign din_3_rsci_biwt = (~ core_wten) & din_3_rsci_oswt;
  assign din_3_rsci_biwt_pff = core_wen & din_3_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1_din_2_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1_din_2_rsc_wait_dp (
  clk, rst, din_2_rsci_douta_d, din_2_rsci_douta_d_mxwt, din_2_rsci_biwt, din_2_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_2_rsci_douta_d;
  output [15:0] din_2_rsci_douta_d_mxwt;
  input din_2_rsci_biwt;
  input din_2_rsci_bdwt;


  // Interconnect Declarations
  reg din_2_rsci_bcwt;
  reg [15:0] din_2_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_2_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_2_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_2_rsci_douta_d[15:0]),
      din_2_rsci_douta_d_bfwt_15_0, din_2_rsci_bcwt);
  assign din_2_rsci_douta_d_mxwt = din_2_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_2_rsci_bcwt <= 1'b0;
      din_2_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_2_rsci_bcwt <= ~((~(din_2_rsci_bcwt | din_2_rsci_biwt)) | din_2_rsci_bdwt);
      din_2_rsci_douta_d_bfwt_15_0 <= din_2_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1_din_2_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1_din_2_rsc_wait_ctrl (
  core_wen, core_wten, din_2_rsci_oswt, din_2_rsci_biwt, din_2_rsci_bdwt, din_2_rsci_biwt_pff,
      din_2_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_2_rsci_oswt;
  output din_2_rsci_biwt;
  output din_2_rsci_bdwt;
  output din_2_rsci_biwt_pff;
  input din_2_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_2_rsci_bdwt = din_2_rsci_oswt & core_wen;
  assign din_2_rsci_biwt = (~ core_wten) & din_2_rsci_oswt;
  assign din_2_rsci_biwt_pff = core_wen & din_2_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1_din_1_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1_din_1_rsc_wait_dp (
  clk, rst, din_1_rsci_douta_d, din_1_rsci_douta_d_mxwt, din_1_rsci_biwt, din_1_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_1_rsci_douta_d;
  output [15:0] din_1_rsci_douta_d_mxwt;
  input din_1_rsci_biwt;
  input din_1_rsci_bdwt;


  // Interconnect Declarations
  reg din_1_rsci_bcwt;
  reg [15:0] din_1_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_1_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_1_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_1_rsci_douta_d[15:0]),
      din_1_rsci_douta_d_bfwt_15_0, din_1_rsci_bcwt);
  assign din_1_rsci_douta_d_mxwt = din_1_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_1_rsci_bcwt <= 1'b0;
      din_1_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_1_rsci_bcwt <= ~((~(din_1_rsci_bcwt | din_1_rsci_biwt)) | din_1_rsci_bdwt);
      din_1_rsci_douta_d_bfwt_15_0 <= din_1_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1_din_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1_din_1_rsc_wait_ctrl (
  core_wen, core_wten, din_1_rsci_oswt, din_1_rsci_biwt, din_1_rsci_bdwt, din_1_rsci_biwt_pff,
      din_1_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_1_rsci_oswt;
  output din_1_rsci_biwt;
  output din_1_rsci_bdwt;
  output din_1_rsci_biwt_pff;
  input din_1_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_1_rsci_bdwt = din_1_rsci_oswt & core_wen;
  assign din_1_rsci_biwt = (~ core_wten) & din_1_rsci_oswt;
  assign din_1_rsci_biwt_pff = core_wen & din_1_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1_din_0_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1_din_0_rsc_wait_dp (
  clk, rst, din_0_rsci_douta_d, din_0_rsci_douta_d_mxwt, din_0_rsci_biwt, din_0_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_0_rsci_douta_d;
  output [15:0] din_0_rsci_douta_d_mxwt;
  input din_0_rsci_biwt;
  input din_0_rsci_bdwt;


  // Interconnect Declarations
  reg din_0_rsci_bcwt;
  reg [15:0] din_0_rsci_douta_d_bfwt_15_0;
  wire [15:0] din_0_rsci_douta_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign din_0_rsci_douta_d_mxwt_opt_15_0 = MUX_v_16_2_2((din_0_rsci_douta_d[15:0]),
      din_0_rsci_douta_d_bfwt_15_0, din_0_rsci_bcwt);
  assign din_0_rsci_douta_d_mxwt = din_0_rsci_douta_d_mxwt_opt_15_0;
  always @(posedge clk) begin
    if ( rst ) begin
      din_0_rsci_bcwt <= 1'b0;
      din_0_rsci_douta_d_bfwt_15_0 <= 16'b0;
    end
    else begin
      din_0_rsci_bcwt <= ~((~(din_0_rsci_bcwt | din_0_rsci_biwt)) | din_0_rsci_bdwt);
      din_0_rsci_douta_d_bfwt_15_0 <= din_0_rsci_douta_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1_din_0_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1_din_0_rsc_wait_ctrl (
  core_wen, din_0_rsci_oswt, core_wten, din_0_rsci_biwt, din_0_rsci_bdwt, din_0_rsci_biwt_pff,
      din_0_rsci_oswt_pff
);
  input core_wen;
  input din_0_rsci_oswt;
  input core_wten;
  output din_0_rsci_biwt;
  output din_0_rsci_bdwt;
  output din_0_rsci_biwt_pff;
  input din_0_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_0_rsci_bdwt = din_0_rsci_oswt & core_wen;
  assign din_0_rsci_biwt = (~ core_wten) & din_0_rsci_oswt;
  assign din_0_rsci_biwt_pff = core_wen & din_0_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffepBGdfem_cns_bctl
// ------------------------------------------------------------------


module double_buffepBGdfem_cns_bctl (
  clk, rst, din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst, dout_rsc_csa_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst,
      dout_rsc_csb_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst, dout_rsc_addra_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst,
      dout_rsc_addrb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst, dout_rsc_dinb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst,
      dout_rsc_douta_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst, dout_rsc_req_vz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst,
      din_rsc_csa_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst, din_rsc_csb_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst,
      din_rsc_addra_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst, din_rsc_addrb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst,
      din_rsc_dinb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst, din_rsc_douta_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst,
      din_rsc_req_vz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst, dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst,
      din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud, dout_rsc_rls_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud,
      din_rsc_rls_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud, dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud,
      shr_mem_cns_S0, shr_mem_cns_R0, shr_mem_cns_S1, shr_mem_cns_R1, shr_mem_cns_addra_shi0,
      shr_mem_cns_addra_shi1, shr_mem_cns_addrb_shi0, shr_mem_cns_addrb_shi1, shr_mem_cns_csa_n_shi0,
      shr_mem_cns_csa_n_shi1, shr_mem_cns_csb_n_shi0, shr_mem_cns_csb_n_shi1, shr_mem_cns_dinb_shi0,
      shr_mem_cns_dinb_shi1, shr_mem_cns_douta_sho0, shr_mem_cns_douta_sho1, shr_mem_cns_S1_pff,
      shr_mem_cns_S0_pff
);
  input clk;
  input rst;
  output din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  input dout_rsc_csa_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  input dout_rsc_csb_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  input [6:0] dout_rsc_addra_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  input [6:0] dout_rsc_addrb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  input [63:0] dout_rsc_dinb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  output [63:0] dout_rsc_douta_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  output dout_rsc_req_vz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  input din_rsc_csa_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  input din_rsc_csb_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  input [6:0] din_rsc_addra_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  input [6:0] din_rsc_addrb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  input [63:0] din_rsc_dinb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  output [63:0] din_rsc_douta_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  output din_rsc_req_vz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  output dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  input din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud;
  input dout_rsc_rls_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud;
  input din_rsc_rls_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud;
  input dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud;
  output shr_mem_cns_S0;
  input shr_mem_cns_R0;
  output shr_mem_cns_S1;
  input shr_mem_cns_R1;
  output [6:0] shr_mem_cns_addra_shi0;
  output [6:0] shr_mem_cns_addra_shi1;
  output [6:0] shr_mem_cns_addrb_shi0;
  output [6:0] shr_mem_cns_addrb_shi1;
  output shr_mem_cns_csa_n_shi0;
  output shr_mem_cns_csa_n_shi1;
  output shr_mem_cns_csb_n_shi0;
  output shr_mem_cns_csb_n_shi1;
  output [63:0] shr_mem_cns_dinb_shi0;
  output [63:0] shr_mem_cns_dinb_shi1;
  input [63:0] shr_mem_cns_douta_sho0;
  input [63:0] shr_mem_cns_douta_sho1;
  output shr_mem_cns_S1_pff;
  output shr_mem_cns_S0_pff;


  // Interconnect Declarations
  wire shr_mem_cns_PC0;
  reg shr_mem_cns_ppidx;
  reg [1:0] shr_mem_cns_ppown;
  wire shr_mem_cns_PC1;
  reg shr_mem_cns_ppidx_1;
  reg [1:0] shr_mem_cns_ppown_1;
  wire [6:0] shr_mem_shr_mem_mux_3_cse_pff;
  wire shr_mem_and_3_cse_pff;
  wire [1:0] shr_mem_acc_1_rmff;
  wire [3:0] nl_shr_mem_acc_1_rmff;
  wire shr_mem_xor_1_rmff;
  wire shr_mem_shr_mem_shr_mem_nand_cse_pff;
  wire [1:0] shr_mem_acc_rmff;
  wire [3:0] nl_shr_mem_acc_rmff;
  wire shr_mem_xor_rmff;
  wire [6:0] shr_mem_shr_mem_mux_2_cse_pff;
  wire shr_mem_and_5_cse_pff;
  wire shr_mem_shr_mem_shr_mem_nand_1_cse_pff;

  wire[0:0] shr_mem_mux_6_nl;
  wire[0:0] shr_mem_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst = din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud;
  assign dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst = dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud;
  assign dout_rsc_req_vz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst = shr_mem_cns_R0;
  assign din_rsc_req_vz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst = shr_mem_cns_R1;
  assign shr_mem_xor_rmff = shr_mem_cns_ppidx ^ shr_mem_cns_PC0;
  assign nl_shr_mem_acc_rmff = shr_mem_cns_ppown + conv_u2u_1_2(shr_mem_cns_PC0)
      + conv_s2u_1_2(shr_mem_cns_PC1);
  assign shr_mem_acc_rmff = nl_shr_mem_acc_rmff[1:0];
  assign shr_mem_cns_PC0 = shr_mem_cns_S0 & dout_rsc_rls_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud;
  assign shr_mem_xor_1_rmff = shr_mem_cns_ppidx_1 ^ shr_mem_cns_PC1;
  assign nl_shr_mem_acc_1_rmff = shr_mem_cns_ppown_1 + conv_u2u_1_2(shr_mem_cns_PC1)
      + conv_s2u_1_2(shr_mem_cns_PC0);
  assign shr_mem_acc_1_rmff = nl_shr_mem_acc_1_rmff[1:0];
  assign shr_mem_cns_PC1 = shr_mem_cns_S1 & din_rsc_rls_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud;
  assign dout_rsc_douta_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst = MUX_v_64_2_2(shr_mem_cns_douta_sho0,
      shr_mem_cns_douta_sho1, shr_mem_cns_ppidx);
  assign din_rsc_douta_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst = MUX_v_64_2_2(shr_mem_cns_douta_sho0,
      shr_mem_cns_douta_sho1, shr_mem_cns_ppidx_1);
  assign shr_mem_cns_addra_shi0 = shr_mem_shr_mem_mux_3_cse_pff;
  assign shr_mem_cns_S1 = (shr_mem_cns_ppown_1!=2'b00);
  assign shr_mem_cns_S1_pff = (shr_mem_acc_1_rmff!=2'b00);
  assign shr_mem_and_3_cse_pff = shr_mem_cns_S1_pff & (~ shr_mem_xor_1_rmff);
  assign shr_mem_shr_mem_mux_3_cse_pff = MUX_v_7_2_2(dout_rsc_addrb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst,
      din_rsc_addrb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst, shr_mem_and_3_cse_pff);
  assign shr_mem_cns_addrb_shi0 = shr_mem_shr_mem_mux_3_cse_pff;
  assign shr_mem_cns_csa_n_shi0 = shr_mem_shr_mem_shr_mem_nand_cse_pff;
  assign shr_mem_cns_S0 = ~((shr_mem_cns_ppown==2'b10));
  assign shr_mem_cns_S0_pff = ~((shr_mem_acc_rmff==2'b10));
  assign shr_mem_mux_6_nl = MUX_s_1_2_2(dout_rsc_csb_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst,
      din_rsc_csb_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst, shr_mem_and_3_cse_pff);
  assign shr_mem_shr_mem_shr_mem_nand_cse_pff = (shr_mem_mux_6_nl) | (~((shr_mem_cns_S0_pff
      & (~ shr_mem_xor_rmff)) | shr_mem_and_3_cse_pff));
  assign shr_mem_cns_csb_n_shi0 = shr_mem_shr_mem_shr_mem_nand_cse_pff;
  assign shr_mem_cns_dinb_shi0 = MUX_v_64_2_2(dout_rsc_dinb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst,
      din_rsc_dinb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst, shr_mem_and_3_cse_pff);
  assign shr_mem_cns_addra_shi1 = shr_mem_shr_mem_mux_2_cse_pff;
  assign shr_mem_and_5_cse_pff = shr_mem_cns_S1_pff & shr_mem_xor_1_rmff;
  assign shr_mem_shr_mem_mux_2_cse_pff = MUX_v_7_2_2(dout_rsc_addrb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst,
      din_rsc_addrb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst, shr_mem_and_5_cse_pff);
  assign shr_mem_cns_addrb_shi1 = shr_mem_shr_mem_mux_2_cse_pff;
  assign shr_mem_cns_csa_n_shi1 = shr_mem_shr_mem_shr_mem_nand_1_cse_pff;
  assign shr_mem_mux_7_nl = MUX_s_1_2_2(dout_rsc_csb_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst,
      din_rsc_csb_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst, shr_mem_and_5_cse_pff);
  assign shr_mem_shr_mem_shr_mem_nand_1_cse_pff = (shr_mem_mux_7_nl) | (~((shr_mem_cns_S0_pff
      & shr_mem_xor_rmff) | shr_mem_and_5_cse_pff));
  assign shr_mem_cns_csb_n_shi1 = shr_mem_shr_mem_shr_mem_nand_1_cse_pff;
  assign shr_mem_cns_dinb_shi1 = MUX_v_64_2_2(dout_rsc_dinb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst,
      din_rsc_dinb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst, shr_mem_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      shr_mem_cns_ppidx <= 1'b0;
      shr_mem_cns_ppown <= 2'b0;
      shr_mem_cns_ppidx_1 <= 1'b0;
      shr_mem_cns_ppown_1 <= 2'b0;
    end
    else begin
      shr_mem_cns_ppidx <= shr_mem_xor_rmff;
      shr_mem_cns_ppown <= shr_mem_acc_rmff;
      shr_mem_cns_ppidx_1 <= shr_mem_xor_1_rmff;
      shr_mem_cns_ppown_1 <= shr_mem_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    unreg_hier_33
// ------------------------------------------------------------------


module unreg_hier_33 (
  in_0, out_0
);
  input in_0;
  output out_0;



  // Interconnect Declarations for Component Instantiations 
  assign out_0 = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_96_n1073741823_0_0_0_36_64_128_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_96_n1073741823_0_0_0_36_64_128_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_and_nl;
  wire dout_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_and_nl);
  assign dout_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_staller
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_staller (
  clk, rst, core_wen, din_rsci_wen_comp, core_wten, dout_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  input din_rsci_wen_comp;
  output core_wten;
  input dout_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = din_rsci_wen_comp & dout_rsc_req_obj_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj_dout_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj_dout_rsc_req_wait_dp
    (
  clk, rst, dout_rsc_req_obj_oswt, dout_rsc_req_obj_wen_comp, dout_rsc_req_obj_biwt,
      dout_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_rsc_req_obj_oswt;
  output dout_rsc_req_obj_wen_comp;
  input dout_rsc_req_obj_biwt;
  input dout_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_req_obj_wen_comp = (~ dout_rsc_req_obj_oswt) | dout_rsc_req_obj_biwt
      | dout_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_rsc_req_obj_bcwt <= ~((~(dout_rsc_req_obj_bcwt | dout_rsc_req_obj_biwt))
          | dout_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_rsc_req_obj_oswt, dout_rsc_req_obj_vd, dout_rsc_req_obj_biwt,
      dout_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_rsc_req_obj_oswt;
  input dout_rsc_req_obj_vd;
  output dout_rsc_req_obj_biwt;
  output dout_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_rsc_req_obj_pdswt0;
  reg dout_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_req_obj_pdswt0 = (~ core_wten) & dout_rsc_req_obj_oswt;
  assign dout_rsc_req_obj_biwt = (dout_rsc_req_obj_pdswt0 | dout_rsc_req_obj_icwt)
      & dout_rsc_req_obj_vd;
  assign dout_rsc_req_obj_bdwt = dout_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_rsc_req_obj_icwt <= ~((~(dout_rsc_req_obj_icwt | dout_rsc_req_obj_pdswt0))
          | dout_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
    (
  core_wten, dout_rsc_rls_obj_iswt0, dout_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_rsc_rls_obj_iswt0;
  output dout_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_rls_obj_ld_core_sct = dout_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_dout_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_dout_rsc_wait_ctrl (
  dout_rsci_addra_d_core_sct_pff, dout_rsci_iswt0_pff, core_wten_pff
);
  output dout_rsci_addra_d_core_sct_pff;
  input dout_rsci_iswt0_pff;
  input core_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_addra_d_core_sct_pff = dout_rsci_iswt0_pff & (~ core_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci_din_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci_din_wait_dp (
  clk, rst, din_rsci_oswt, din_rsci_wen_comp, din_rsci_d_mxwt, din_rsci_biwt, din_rsci_bdwt,
      din_rsci_d
);
  input clk;
  input rst;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [63:0] din_rsci_d_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  input [63:0] din_rsci_d;


  // Interconnect Declarations
  reg din_rsci_bcwt;
  reg [63:0] din_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_wen_comp = (~ din_rsci_oswt) | din_rsci_biwt | din_rsci_bcwt;
  assign din_rsci_d_mxwt = MUX_v_64_2_2(din_rsci_d, din_rsci_d_bfwt, din_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsci_bcwt <= 1'b0;
      din_rsci_d_bfwt <= 64'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
      din_rsci_d_bfwt <= din_rsci_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci_din_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci_din_wait_ctrl (
  clk, rst, core_wen, din_rsci_oswt, core_wten, din_rsci_biwt, din_rsci_bdwt, din_rsci_ld_core_sct,
      din_rsci_vd
);
  input clk;
  input rst;
  input core_wen;
  input din_rsci_oswt;
  input core_wten;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  output din_rsci_ld_core_sct;
  input din_rsci_vd;


  // Interconnect Declarations
  wire din_rsci_ogwt;
  wire din_rsci_pdswt0;
  reg din_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_pdswt0 = (~ core_wten) & din_rsci_oswt;
  assign din_rsci_biwt = din_rsci_ogwt & din_rsci_vd;
  assign din_rsci_ogwt = din_rsci_pdswt0 | din_rsci_icwt;
  assign din_rsci_bdwt = din_rsci_oswt & core_wen;
  assign din_rsci_ld_core_sct = din_rsci_oswt & din_rsci_ogwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsci_icwt <= 1'b0;
    end
    else begin
      din_rsci_icwt <= ~((~(din_rsci_icwt | din_rsci_pdswt0)) | din_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_98_n1073741823_0_0_0_36_64_128_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_98_n1073741823_0_0_0_36_64_128_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [6:0] addrb;
  output [6:0] addra;
  output csb_n;
  output csa_n;
  input [6:0] addra_d;
  input [6:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_and_nl;
  wire din_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_and_nl);
  assign din_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_staller
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_staller (
  clk, rst, core_wen, core_wten, dout_rsci_wen_comp, din_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input dout_rsci_wen_comp;
  input din_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = dout_rsci_wen_comp & din_rsc_req_obj_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj_din_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj_din_rsc_req_wait_dp
    (
  clk, rst, din_rsc_req_obj_oswt, din_rsc_req_obj_wen_comp, din_rsc_req_obj_biwt,
      din_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_rsc_req_obj_oswt;
  output din_rsc_req_obj_wen_comp;
  input din_rsc_req_obj_biwt;
  input din_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_req_obj_wen_comp = (~ din_rsc_req_obj_oswt) | din_rsc_req_obj_biwt
      | din_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_rsc_req_obj_bcwt <= ~((~(din_rsc_req_obj_bcwt | din_rsc_req_obj_biwt))
          | din_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj_din_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj_din_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_rsc_req_obj_oswt, din_rsc_req_obj_vd, din_rsc_req_obj_biwt,
      din_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_rsc_req_obj_oswt;
  input din_rsc_req_obj_vd;
  output din_rsc_req_obj_biwt;
  output din_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_rsc_req_obj_pdswt0;
  reg din_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_req_obj_pdswt0 = (~ core_wten) & din_rsc_req_obj_oswt;
  assign din_rsc_req_obj_biwt = (din_rsc_req_obj_pdswt0 | din_rsc_req_obj_icwt) &
      din_rsc_req_obj_vd;
  assign din_rsc_req_obj_bdwt = din_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_rsc_req_obj_icwt <= ~((~(din_rsc_req_obj_icwt | din_rsc_req_obj_pdswt0))
          | din_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
    (
  core_wten, din_rsc_rls_obj_iswt0, din_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_rsc_rls_obj_iswt0;
  output din_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_rls_obj_ld_core_sct = din_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci_dout_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci_dout_wait_dp (
  clk, rst, dout_rsci_oswt, dout_rsci_wen_comp, dout_rsci_biwt, dout_rsci_bdwt
);
  input clk;
  input rst;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input dout_rsci_biwt;
  input dout_rsci_bdwt;


  // Interconnect Declarations
  reg dout_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_wen_comp = (~ dout_rsci_oswt) | dout_rsci_biwt | dout_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_bcwt <= 1'b0;
    end
    else begin
      dout_rsci_bcwt <= ~((~(dout_rsci_bcwt | dout_rsci_biwt)) | dout_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci_dout_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci_dout_wait_ctrl (
  clk, rst, core_wen, core_wten, dout_rsci_oswt, dout_rsci_biwt, dout_rsci_bdwt,
      dout_rsci_ld_core_sct, dout_rsci_vd
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_rsci_oswt;
  output dout_rsci_biwt;
  output dout_rsci_bdwt;
  output dout_rsci_ld_core_sct;
  input dout_rsci_vd;


  // Interconnect Declarations
  wire dout_rsci_ogwt;
  wire dout_rsci_pdswt0;
  reg dout_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_pdswt0 = (~ core_wten) & dout_rsci_oswt;
  assign dout_rsci_biwt = dout_rsci_ogwt & dout_rsci_vd;
  assign dout_rsci_ogwt = dout_rsci_pdswt0 | dout_rsci_icwt;
  assign dout_rsci_bdwt = dout_rsci_oswt & core_wen;
  assign dout_rsci_ld_core_sct = dout_rsci_oswt & dout_rsci_ogwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_icwt <= 1'b0;
    end
    else begin
      dout_rsci_icwt <= ~((~(dout_rsci_icwt | dout_rsci_pdswt0)) | dout_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_dp (
  clk, rst, din_rsci_addra_d, din_rsci_addrb_d, din_rsci_douta_d, din_rsci_addra_d_core,
      din_rsci_addrb_d_core, din_rsci_douta_d_mxwt, din_rsci_biwt, din_rsci_bdwt,
      din_rsci_biwt_pff
);
  input clk;
  input rst;
  output [6:0] din_rsci_addra_d;
  output [6:0] din_rsci_addrb_d;
  input [63:0] din_rsci_douta_d;
  input [6:0] din_rsci_addra_d_core;
  input [6:0] din_rsci_addrb_d_core;
  output [63:0] din_rsci_douta_d_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  input din_rsci_biwt_pff;


  // Interconnect Declarations
  reg din_rsci_bcwt;
  reg [63:0] din_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_douta_d_mxwt = MUX_v_64_2_2(din_rsci_douta_d, din_rsci_douta_d_bfwt,
      din_rsci_bcwt);
  assign din_rsci_addra_d = {(~ din_rsci_biwt_pff) , (din_rsci_addra_d_core[5:0])};
  assign din_rsci_addrb_d = {(~ din_rsci_biwt_pff) , (din_rsci_addrb_d_core[5:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsci_bcwt <= 1'b0;
      din_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
      din_rsci_douta_d_bfwt <= din_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_ctrl (
  core_wen, din_rsci_oswt, core_wten, din_rsci_biwt, din_rsci_bdwt, din_rsci_biwt_pff,
      din_rsci_oswt_pff
);
  input core_wen;
  input din_rsci_oswt;
  input core_wten;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  output din_rsci_biwt_pff;
  input din_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_bdwt = din_rsci_oswt & core_wen;
  assign din_rsci_biwt = (~ core_wten) & din_rsci_oswt;
  assign din_rsci_biwt_pff = core_wen & din_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core_staller
// ------------------------------------------------------------------


module systolic_array_core_staller (
  clk, rst, core_wen, input_rsci_wen_comp, core_wten, weight_rsci_wen_comp, output_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  input input_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input weight_rsci_wen_comp;
  input output_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = input_rsci_wen_comp & weight_rsci_wen_comp & output_rsci_wen_comp;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core_output_rsci_output_wait_dp
// ------------------------------------------------------------------


module systolic_array_core_output_rsci_output_wait_dp (
  clk, rst, output_rsci_oswt, output_rsci_wen_comp, output_rsci_biwt, output_rsci_bdwt
);
  input clk;
  input rst;
  input output_rsci_oswt;
  output output_rsci_wen_comp;
  input output_rsci_biwt;
  input output_rsci_bdwt;


  // Interconnect Declarations
  reg output_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_rsci_wen_comp = (~ output_rsci_oswt) | output_rsci_biwt | output_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_bcwt <= 1'b0;
    end
    else begin
      output_rsci_bcwt <= ~((~(output_rsci_bcwt | output_rsci_biwt)) | output_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core_output_rsci_output_wait_ctrl
// ------------------------------------------------------------------


module systolic_array_core_output_rsci_output_wait_ctrl (
  clk, rst, core_wen, core_wten, output_rsci_oswt, output_rsci_biwt, output_rsci_bdwt,
      output_rsci_ld_core_sct, output_rsci_vd
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input output_rsci_oswt;
  output output_rsci_biwt;
  output output_rsci_bdwt;
  output output_rsci_ld_core_sct;
  input output_rsci_vd;


  // Interconnect Declarations
  wire output_rsci_ogwt;
  wire output_rsci_pdswt0;
  reg output_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_rsci_pdswt0 = (~ core_wten) & output_rsci_oswt;
  assign output_rsci_biwt = output_rsci_ogwt & output_rsci_vd;
  assign output_rsci_ogwt = output_rsci_pdswt0 | output_rsci_icwt;
  assign output_rsci_bdwt = output_rsci_oswt & core_wen;
  assign output_rsci_ld_core_sct = output_rsci_oswt & output_rsci_ogwt;
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_icwt <= 1'b0;
    end
    else begin
      output_rsci_icwt <= ~((~(output_rsci_icwt | output_rsci_pdswt0)) | output_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core_weight_rsci_weight_wait_dp
// ------------------------------------------------------------------


module systolic_array_core_weight_rsci_weight_wait_dp (
  clk, rst, weight_rsci_oswt, weight_rsci_wen_comp, weight_rsci_d_mxwt, weight_rsci_biwt,
      weight_rsci_bdwt, weight_rsci_d
);
  input clk;
  input rst;
  input weight_rsci_oswt;
  output weight_rsci_wen_comp;
  output [31:0] weight_rsci_d_mxwt;
  input weight_rsci_biwt;
  input weight_rsci_bdwt;
  input [63:0] weight_rsci_d;


  // Interconnect Declarations
  reg weight_rsci_bcwt;
  reg [15:0] reg_weight_rsci_d_bfwt_tmp;
  reg [15:0] reg_weight_rsci_d_bfwt_tmp_17;
  wire [15:0] weight_rsci_d_mxwt_opt_47_32;
  wire [15:0] weight_rsci_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign weight_rsci_wen_comp = (~ weight_rsci_oswt) | weight_rsci_biwt | weight_rsci_bcwt;
  assign weight_rsci_d_mxwt_opt_47_32 = MUX_v_16_2_2((weight_rsci_d[47:32]), reg_weight_rsci_d_bfwt_tmp,
      weight_rsci_bcwt);
  assign weight_rsci_d_mxwt_opt_15_0 = MUX_v_16_2_2((weight_rsci_d[15:0]), reg_weight_rsci_d_bfwt_tmp_17,
      weight_rsci_bcwt);
  assign weight_rsci_d_mxwt = {weight_rsci_d_mxwt_opt_47_32 , weight_rsci_d_mxwt_opt_15_0};
  always @(posedge clk) begin
    if ( rst ) begin
      weight_rsci_bcwt <= 1'b0;
      reg_weight_rsci_d_bfwt_tmp <= 16'b0;
      reg_weight_rsci_d_bfwt_tmp_17 <= 16'b0;
    end
    else begin
      weight_rsci_bcwt <= ~((~(weight_rsci_bcwt | weight_rsci_biwt)) | weight_rsci_bdwt);
      reg_weight_rsci_d_bfwt_tmp <= weight_rsci_d_mxwt_opt_47_32;
      reg_weight_rsci_d_bfwt_tmp_17 <= weight_rsci_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core_weight_rsci_weight_wait_ctrl
// ------------------------------------------------------------------


module systolic_array_core_weight_rsci_weight_wait_ctrl (
  clk, rst, core_wen, core_wten, weight_rsci_oswt, weight_rsci_biwt, weight_rsci_bdwt,
      weight_rsci_ld_core_sct, weight_rsci_vd
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input weight_rsci_oswt;
  output weight_rsci_biwt;
  output weight_rsci_bdwt;
  output weight_rsci_ld_core_sct;
  input weight_rsci_vd;


  // Interconnect Declarations
  wire weight_rsci_ogwt;
  wire weight_rsci_pdswt0;
  reg weight_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign weight_rsci_pdswt0 = (~ core_wten) & weight_rsci_oswt;
  assign weight_rsci_biwt = weight_rsci_ogwt & weight_rsci_vd;
  assign weight_rsci_ogwt = weight_rsci_pdswt0 | weight_rsci_icwt;
  assign weight_rsci_bdwt = weight_rsci_oswt & core_wen;
  assign weight_rsci_ld_core_sct = weight_rsci_oswt & weight_rsci_ogwt;
  always @(posedge clk) begin
    if ( rst ) begin
      weight_rsci_icwt <= 1'b0;
    end
    else begin
      weight_rsci_icwt <= ~((~(weight_rsci_icwt | weight_rsci_pdswt0)) | weight_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core_input_rsci_input_wait_dp
// ------------------------------------------------------------------


module systolic_array_core_input_rsci_input_wait_dp (
  clk, rst, input_rsci_oswt, input_rsci_wen_comp, input_rsci_d_mxwt, input_rsci_biwt,
      input_rsci_bdwt, input_rsci_d
);
  input clk;
  input rst;
  input input_rsci_oswt;
  output input_rsci_wen_comp;
  output [255:0] input_rsci_d_mxwt;
  input input_rsci_biwt;
  input input_rsci_bdwt;
  input [511:0] input_rsci_d;


  // Interconnect Declarations
  reg input_rsci_bcwt;
  reg [15:0] reg_input_rsci_d_bfwt_tmp;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_17;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_34;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_51;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_68;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_85;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_102;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_119;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_136;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_153;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_170;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_187;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_204;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_221;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_238;
  reg [15:0] reg_input_rsci_d_bfwt_tmp_255;
  wire [15:0] input_rsci_d_mxwt_opt_495_480;
  wire [15:0] input_rsci_d_mxwt_opt_463_448;
  wire [15:0] input_rsci_d_mxwt_opt_431_416;
  wire [15:0] input_rsci_d_mxwt_opt_399_384;
  wire [15:0] input_rsci_d_mxwt_opt_367_352;
  wire [15:0] input_rsci_d_mxwt_opt_335_320;
  wire [15:0] input_rsci_d_mxwt_opt_303_288;
  wire [15:0] input_rsci_d_mxwt_opt_271_256;
  wire [15:0] input_rsci_d_mxwt_opt_239_224;
  wire [15:0] input_rsci_d_mxwt_opt_207_192;
  wire [15:0] input_rsci_d_mxwt_opt_175_160;
  wire [15:0] input_rsci_d_mxwt_opt_143_128;
  wire [15:0] input_rsci_d_mxwt_opt_111_96;
  wire [15:0] input_rsci_d_mxwt_opt_79_64;
  wire [15:0] input_rsci_d_mxwt_opt_47_32;
  wire [15:0] input_rsci_d_mxwt_opt_15_0;


  // Interconnect Declarations for Component Instantiations 
  assign input_rsci_wen_comp = (~ input_rsci_oswt) | input_rsci_biwt | input_rsci_bcwt;
  assign input_rsci_d_mxwt_opt_495_480 = MUX_v_16_2_2((input_rsci_d[495:480]), reg_input_rsci_d_bfwt_tmp,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_463_448 = MUX_v_16_2_2((input_rsci_d[463:448]), reg_input_rsci_d_bfwt_tmp_17,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_431_416 = MUX_v_16_2_2((input_rsci_d[431:416]), reg_input_rsci_d_bfwt_tmp_34,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_399_384 = MUX_v_16_2_2((input_rsci_d[399:384]), reg_input_rsci_d_bfwt_tmp_51,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_367_352 = MUX_v_16_2_2((input_rsci_d[367:352]), reg_input_rsci_d_bfwt_tmp_68,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_335_320 = MUX_v_16_2_2((input_rsci_d[335:320]), reg_input_rsci_d_bfwt_tmp_85,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_303_288 = MUX_v_16_2_2((input_rsci_d[303:288]), reg_input_rsci_d_bfwt_tmp_102,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_271_256 = MUX_v_16_2_2((input_rsci_d[271:256]), reg_input_rsci_d_bfwt_tmp_119,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_239_224 = MUX_v_16_2_2((input_rsci_d[239:224]), reg_input_rsci_d_bfwt_tmp_136,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_207_192 = MUX_v_16_2_2((input_rsci_d[207:192]), reg_input_rsci_d_bfwt_tmp_153,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_175_160 = MUX_v_16_2_2((input_rsci_d[175:160]), reg_input_rsci_d_bfwt_tmp_170,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_143_128 = MUX_v_16_2_2((input_rsci_d[143:128]), reg_input_rsci_d_bfwt_tmp_187,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_111_96 = MUX_v_16_2_2((input_rsci_d[111:96]), reg_input_rsci_d_bfwt_tmp_204,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_79_64 = MUX_v_16_2_2((input_rsci_d[79:64]), reg_input_rsci_d_bfwt_tmp_221,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_47_32 = MUX_v_16_2_2((input_rsci_d[47:32]), reg_input_rsci_d_bfwt_tmp_238,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt_opt_15_0 = MUX_v_16_2_2((input_rsci_d[15:0]), reg_input_rsci_d_bfwt_tmp_255,
      input_rsci_bcwt);
  assign input_rsci_d_mxwt = {input_rsci_d_mxwt_opt_495_480 , input_rsci_d_mxwt_opt_463_448
      , input_rsci_d_mxwt_opt_431_416 , input_rsci_d_mxwt_opt_399_384 , input_rsci_d_mxwt_opt_367_352
      , input_rsci_d_mxwt_opt_335_320 , input_rsci_d_mxwt_opt_303_288 , input_rsci_d_mxwt_opt_271_256
      , input_rsci_d_mxwt_opt_239_224 , input_rsci_d_mxwt_opt_207_192 , input_rsci_d_mxwt_opt_175_160
      , input_rsci_d_mxwt_opt_143_128 , input_rsci_d_mxwt_opt_111_96 , input_rsci_d_mxwt_opt_79_64
      , input_rsci_d_mxwt_opt_47_32 , input_rsci_d_mxwt_opt_15_0};
  always @(posedge clk) begin
    if ( rst ) begin
      input_rsci_bcwt <= 1'b0;
      reg_input_rsci_d_bfwt_tmp <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_17 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_34 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_51 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_68 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_85 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_102 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_119 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_136 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_153 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_170 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_187 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_204 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_221 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_238 <= 16'b0;
      reg_input_rsci_d_bfwt_tmp_255 <= 16'b0;
    end
    else begin
      input_rsci_bcwt <= ~((~(input_rsci_bcwt | input_rsci_biwt)) | input_rsci_bdwt);
      reg_input_rsci_d_bfwt_tmp <= input_rsci_d_mxwt_opt_495_480;
      reg_input_rsci_d_bfwt_tmp_17 <= input_rsci_d_mxwt_opt_463_448;
      reg_input_rsci_d_bfwt_tmp_34 <= input_rsci_d_mxwt_opt_431_416;
      reg_input_rsci_d_bfwt_tmp_51 <= input_rsci_d_mxwt_opt_399_384;
      reg_input_rsci_d_bfwt_tmp_68 <= input_rsci_d_mxwt_opt_367_352;
      reg_input_rsci_d_bfwt_tmp_85 <= input_rsci_d_mxwt_opt_335_320;
      reg_input_rsci_d_bfwt_tmp_102 <= input_rsci_d_mxwt_opt_303_288;
      reg_input_rsci_d_bfwt_tmp_119 <= input_rsci_d_mxwt_opt_271_256;
      reg_input_rsci_d_bfwt_tmp_136 <= input_rsci_d_mxwt_opt_239_224;
      reg_input_rsci_d_bfwt_tmp_153 <= input_rsci_d_mxwt_opt_207_192;
      reg_input_rsci_d_bfwt_tmp_170 <= input_rsci_d_mxwt_opt_175_160;
      reg_input_rsci_d_bfwt_tmp_187 <= input_rsci_d_mxwt_opt_143_128;
      reg_input_rsci_d_bfwt_tmp_204 <= input_rsci_d_mxwt_opt_111_96;
      reg_input_rsci_d_bfwt_tmp_221 <= input_rsci_d_mxwt_opt_79_64;
      reg_input_rsci_d_bfwt_tmp_238 <= input_rsci_d_mxwt_opt_47_32;
      reg_input_rsci_d_bfwt_tmp_255 <= input_rsci_d_mxwt_opt_15_0;
    end
  end

  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core_input_rsci_input_wait_ctrl
// ------------------------------------------------------------------


module systolic_array_core_input_rsci_input_wait_ctrl (
  clk, rst, core_wen, input_rsci_oswt, core_wten, input_rsci_biwt, input_rsci_bdwt,
      input_rsci_ld_core_sct, input_rsci_vd
);
  input clk;
  input rst;
  input core_wen;
  input input_rsci_oswt;
  input core_wten;
  output input_rsci_biwt;
  output input_rsci_bdwt;
  output input_rsci_ld_core_sct;
  input input_rsci_vd;


  // Interconnect Declarations
  wire input_rsci_ogwt;
  wire input_rsci_pdswt0;
  reg input_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_rsci_pdswt0 = (~ core_wten) & input_rsci_oswt;
  assign input_rsci_biwt = input_rsci_ogwt & input_rsci_vd;
  assign input_rsci_ogwt = input_rsci_pdswt0 | input_rsci_icwt;
  assign input_rsci_bdwt = input_rsci_oswt & core_wen;
  assign input_rsci_ld_core_sct = input_rsci_oswt & input_rsci_ogwt;
  always @(posedge clk) begin
    if ( rst ) begin
      input_rsci_icwt <= 1'b0;
    end
    else begin
      input_rsci_icwt <= ~((~(input_rsci_icwt | input_rsci_pdswt0)) | input_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffefnCNP15_cns_bctl
// ------------------------------------------------------------------


module double_buffefnCNP15_cns_bctl (
  clk, rst, dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_15_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_15_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_15_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_15_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_15_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_15_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_15_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_15_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_15_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_15_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_15_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_15_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_15_cns_S0, shr_mem_15_cns_R0, shr_mem_15_cns_S1, shr_mem_15_cns_R1,
      shr_mem_15_cns_addra_shi0, shr_mem_15_cns_addra_shi1, shr_mem_15_cns_addrb_shi0,
      shr_mem_15_cns_addrb_shi1, shr_mem_15_cns_csa_n_shi0, shr_mem_15_cns_csa_n_shi1,
      shr_mem_15_cns_csb_n_shi0, shr_mem_15_cns_csb_n_shi1, shr_mem_15_cns_dinb_shi0,
      shr_mem_15_cns_dinb_shi1, shr_mem_15_cns_douta_sho0, shr_mem_15_cns_douta_sho1,
      shr_mem_15_cns_S1_pff, din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_15_cns_S0_pff
);
  input clk;
  input rst;
  input dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_15_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_15_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_15_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_15_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_15_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_15_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_15_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_15_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_15_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_15_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_15_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_15_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_15_cns_S0;
  input shr_mem_15_cns_R0;
  output shr_mem_15_cns_S1;
  input shr_mem_15_cns_R1;
  output [7:0] shr_mem_15_cns_addra_shi0;
  output [7:0] shr_mem_15_cns_addra_shi1;
  output [7:0] shr_mem_15_cns_addrb_shi0;
  output [7:0] shr_mem_15_cns_addrb_shi1;
  output shr_mem_15_cns_csa_n_shi0;
  output shr_mem_15_cns_csa_n_shi1;
  output shr_mem_15_cns_csb_n_shi0;
  output shr_mem_15_cns_csb_n_shi1;
  output [63:0] shr_mem_15_cns_dinb_shi0;
  output [63:0] shr_mem_15_cns_dinb_shi1;
  input [63:0] shr_mem_15_cns_douta_sho0;
  input [63:0] shr_mem_15_cns_douta_sho1;
  output shr_mem_15_cns_S1_pff;
  input din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_15_cns_S0_pff;


  // Interconnect Declarations
  reg dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_15_cns_PC0;
  reg shr_mem_15_cns_ppidx;
  reg [1:0] shr_mem_15_cns_ppown;
  wire shr_mem_15_cns_PC1;
  reg shr_mem_15_cns_ppidx_1;
  reg [1:0] shr_mem_15_cns_ppown_1;
  wire [7:0] shr_mem_15_shr_mem_15_mux_3_cse_pff;
  wire shr_mem_15_and_3_cse_pff;
  wire [1:0] shr_mem_15_acc_1_rmff;
  wire [3:0] nl_shr_mem_15_acc_1_rmff;
  wire shr_mem_15_xor_1_rmff;
  wire shr_mem_15_shr_mem_15_or_cse_pff;
  wire [1:0] shr_mem_15_acc_rmff;
  wire [3:0] nl_shr_mem_15_acc_rmff;
  wire shr_mem_15_xor_rmff;
  wire [7:0] shr_mem_15_shr_mem_15_mux_2_cse_pff;
  wire shr_mem_15_and_5_cse_pff;
  wire shr_mem_15_shr_mem_15_or_1_cse_pff;

  wire[0:0] shr_mem_15_mux_6_nl;
  wire[0:0] shr_mem_15_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_15_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_15_cns_R0;
  assign din_15_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_15_cns_R1;
  assign shr_mem_15_xor_rmff = shr_mem_15_cns_ppidx ^ shr_mem_15_cns_PC0;
  assign nl_shr_mem_15_acc_rmff = shr_mem_15_cns_ppown + conv_u2u_1_2(shr_mem_15_cns_PC0)
      + conv_s2u_1_2(shr_mem_15_cns_PC1);
  assign shr_mem_15_acc_rmff = nl_shr_mem_15_acc_rmff[1:0];
  assign shr_mem_15_cns_PC0 = shr_mem_15_cns_S0 & dout_15_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_15_xor_1_rmff = shr_mem_15_cns_ppidx_1 ^ shr_mem_15_cns_PC1;
  assign nl_shr_mem_15_acc_1_rmff = shr_mem_15_cns_ppown_1 + conv_u2u_1_2(shr_mem_15_cns_PC1)
      + conv_s2u_1_2(shr_mem_15_cns_PC0);
  assign shr_mem_15_acc_1_rmff = nl_shr_mem_15_acc_1_rmff[1:0];
  assign shr_mem_15_cns_PC1 = shr_mem_15_cns_S1 & din_15_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_15_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_15_cns_douta_sho0,
      shr_mem_15_cns_douta_sho1, shr_mem_15_cns_ppidx);
  assign din_15_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_15_cns_douta_sho0,
      shr_mem_15_cns_douta_sho1, shr_mem_15_cns_ppidx_1);
  assign shr_mem_15_cns_addra_shi0 = shr_mem_15_shr_mem_15_mux_3_cse_pff;
  assign shr_mem_15_cns_S1 = (shr_mem_15_cns_ppown_1!=2'b00);
  assign shr_mem_15_cns_S1_pff = (shr_mem_15_acc_1_rmff!=2'b00);
  assign shr_mem_15_and_3_cse_pff = shr_mem_15_cns_S1_pff & (~ shr_mem_15_xor_1_rmff);
  assign shr_mem_15_shr_mem_15_mux_3_cse_pff = MUX_v_8_2_2(dout_15_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_15_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_15_and_3_cse_pff);
  assign shr_mem_15_cns_addrb_shi0 = shr_mem_15_shr_mem_15_mux_3_cse_pff;
  assign shr_mem_15_cns_csa_n_shi0 = shr_mem_15_shr_mem_15_or_cse_pff;
  assign din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_15_cns_S0 = ~((shr_mem_15_cns_ppown==2'b10));
  assign shr_mem_15_cns_S0_pff = ~((shr_mem_15_acc_rmff==2'b10));
  assign shr_mem_15_mux_6_nl = MUX_s_1_2_2(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_15_and_3_cse_pff);
  assign shr_mem_15_shr_mem_15_or_cse_pff = (shr_mem_15_mux_6_nl) | (~((shr_mem_15_cns_S0_pff
      & (~ shr_mem_15_xor_rmff)) | shr_mem_15_and_3_cse_pff));
  assign shr_mem_15_cns_csb_n_shi0 = shr_mem_15_shr_mem_15_or_cse_pff;
  assign shr_mem_15_cns_dinb_shi0 = MUX_v_64_2_2(dout_15_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_15_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_15_and_3_cse_pff);
  assign shr_mem_15_cns_addra_shi1 = shr_mem_15_shr_mem_15_mux_2_cse_pff;
  assign shr_mem_15_and_5_cse_pff = shr_mem_15_cns_S1_pff & shr_mem_15_xor_1_rmff;
  assign shr_mem_15_shr_mem_15_mux_2_cse_pff = MUX_v_8_2_2(dout_15_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_15_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_15_and_5_cse_pff);
  assign shr_mem_15_cns_addrb_shi1 = shr_mem_15_shr_mem_15_mux_2_cse_pff;
  assign shr_mem_15_cns_csa_n_shi1 = shr_mem_15_shr_mem_15_or_1_cse_pff;
  assign shr_mem_15_mux_7_nl = MUX_s_1_2_2(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_15_and_5_cse_pff);
  assign shr_mem_15_shr_mem_15_or_1_cse_pff = (shr_mem_15_mux_7_nl) | (~((shr_mem_15_cns_S0_pff
      & shr_mem_15_xor_rmff) | shr_mem_15_and_5_cse_pff));
  assign shr_mem_15_cns_csb_n_shi1 = shr_mem_15_shr_mem_15_or_1_cse_pff;
  assign shr_mem_15_cns_dinb_shi1 = MUX_v_64_2_2(dout_15_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_15_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_15_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_15_cns_ppidx <= 1'b0;
      shr_mem_15_cns_ppown <= 2'b0;
      shr_mem_15_cns_ppidx_1 <= 1'b0;
      shr_mem_15_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_15_cns_ppidx <= shr_mem_15_xor_rmff;
      shr_mem_15_cns_ppown <= shr_mem_15_acc_rmff;
      shr_mem_15_cns_ppidx_1 <= shr_mem_15_xor_1_rmff;
      shr_mem_15_cns_ppown_1 <= shr_mem_15_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffefnCNP14_cns_bctl
// ------------------------------------------------------------------


module double_buffefnCNP14_cns_bctl (
  clk, rst, dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_14_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_14_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_14_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_14_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_14_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_14_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_14_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_14_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_14_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_14_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_14_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_14_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_14_cns_S0, shr_mem_14_cns_R0, shr_mem_14_cns_S1, shr_mem_14_cns_R1,
      shr_mem_14_cns_addra_shi0, shr_mem_14_cns_addra_shi1, shr_mem_14_cns_addrb_shi0,
      shr_mem_14_cns_addrb_shi1, shr_mem_14_cns_csa_n_shi0, shr_mem_14_cns_csa_n_shi1,
      shr_mem_14_cns_csb_n_shi0, shr_mem_14_cns_csb_n_shi1, shr_mem_14_cns_dinb_shi0,
      shr_mem_14_cns_dinb_shi1, shr_mem_14_cns_douta_sho0, shr_mem_14_cns_douta_sho1,
      shr_mem_14_cns_S1_pff, din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_14_cns_S0_pff
);
  input clk;
  input rst;
  input dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_14_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_14_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_14_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_14_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_14_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_14_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_14_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_14_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_14_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_14_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_14_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_14_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_14_cns_S0;
  input shr_mem_14_cns_R0;
  output shr_mem_14_cns_S1;
  input shr_mem_14_cns_R1;
  output [7:0] shr_mem_14_cns_addra_shi0;
  output [7:0] shr_mem_14_cns_addra_shi1;
  output [7:0] shr_mem_14_cns_addrb_shi0;
  output [7:0] shr_mem_14_cns_addrb_shi1;
  output shr_mem_14_cns_csa_n_shi0;
  output shr_mem_14_cns_csa_n_shi1;
  output shr_mem_14_cns_csb_n_shi0;
  output shr_mem_14_cns_csb_n_shi1;
  output [63:0] shr_mem_14_cns_dinb_shi0;
  output [63:0] shr_mem_14_cns_dinb_shi1;
  input [63:0] shr_mem_14_cns_douta_sho0;
  input [63:0] shr_mem_14_cns_douta_sho1;
  output shr_mem_14_cns_S1_pff;
  input din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_14_cns_S0_pff;


  // Interconnect Declarations
  reg dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_14_cns_PC0;
  reg shr_mem_14_cns_ppidx;
  reg [1:0] shr_mem_14_cns_ppown;
  wire shr_mem_14_cns_PC1;
  reg shr_mem_14_cns_ppidx_1;
  reg [1:0] shr_mem_14_cns_ppown_1;
  wire [7:0] shr_mem_14_shr_mem_14_mux_3_cse_pff;
  wire shr_mem_14_and_3_cse_pff;
  wire [1:0] shr_mem_14_acc_1_rmff;
  wire [3:0] nl_shr_mem_14_acc_1_rmff;
  wire shr_mem_14_xor_1_rmff;
  wire shr_mem_14_shr_mem_14_or_cse_pff;
  wire [1:0] shr_mem_14_acc_rmff;
  wire [3:0] nl_shr_mem_14_acc_rmff;
  wire shr_mem_14_xor_rmff;
  wire [7:0] shr_mem_14_shr_mem_14_mux_2_cse_pff;
  wire shr_mem_14_and_5_cse_pff;
  wire shr_mem_14_shr_mem_14_or_1_cse_pff;

  wire[0:0] shr_mem_14_mux_6_nl;
  wire[0:0] shr_mem_14_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_14_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_14_cns_R0;
  assign din_14_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_14_cns_R1;
  assign shr_mem_14_xor_rmff = shr_mem_14_cns_ppidx ^ shr_mem_14_cns_PC0;
  assign nl_shr_mem_14_acc_rmff = shr_mem_14_cns_ppown + conv_u2u_1_2(shr_mem_14_cns_PC0)
      + conv_s2u_1_2(shr_mem_14_cns_PC1);
  assign shr_mem_14_acc_rmff = nl_shr_mem_14_acc_rmff[1:0];
  assign shr_mem_14_cns_PC0 = shr_mem_14_cns_S0 & dout_14_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_14_xor_1_rmff = shr_mem_14_cns_ppidx_1 ^ shr_mem_14_cns_PC1;
  assign nl_shr_mem_14_acc_1_rmff = shr_mem_14_cns_ppown_1 + conv_u2u_1_2(shr_mem_14_cns_PC1)
      + conv_s2u_1_2(shr_mem_14_cns_PC0);
  assign shr_mem_14_acc_1_rmff = nl_shr_mem_14_acc_1_rmff[1:0];
  assign shr_mem_14_cns_PC1 = shr_mem_14_cns_S1 & din_14_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_14_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_14_cns_douta_sho0,
      shr_mem_14_cns_douta_sho1, shr_mem_14_cns_ppidx);
  assign din_14_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_14_cns_douta_sho0,
      shr_mem_14_cns_douta_sho1, shr_mem_14_cns_ppidx_1);
  assign shr_mem_14_cns_addra_shi0 = shr_mem_14_shr_mem_14_mux_3_cse_pff;
  assign shr_mem_14_cns_S1 = (shr_mem_14_cns_ppown_1!=2'b00);
  assign shr_mem_14_cns_S1_pff = (shr_mem_14_acc_1_rmff!=2'b00);
  assign shr_mem_14_and_3_cse_pff = shr_mem_14_cns_S1_pff & (~ shr_mem_14_xor_1_rmff);
  assign shr_mem_14_shr_mem_14_mux_3_cse_pff = MUX_v_8_2_2(dout_14_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_14_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_14_and_3_cse_pff);
  assign shr_mem_14_cns_addrb_shi0 = shr_mem_14_shr_mem_14_mux_3_cse_pff;
  assign shr_mem_14_cns_csa_n_shi0 = shr_mem_14_shr_mem_14_or_cse_pff;
  assign din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_14_cns_S0 = ~((shr_mem_14_cns_ppown==2'b10));
  assign shr_mem_14_cns_S0_pff = ~((shr_mem_14_acc_rmff==2'b10));
  assign shr_mem_14_mux_6_nl = MUX_s_1_2_2(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_14_and_3_cse_pff);
  assign shr_mem_14_shr_mem_14_or_cse_pff = (shr_mem_14_mux_6_nl) | (~((shr_mem_14_cns_S0_pff
      & (~ shr_mem_14_xor_rmff)) | shr_mem_14_and_3_cse_pff));
  assign shr_mem_14_cns_csb_n_shi0 = shr_mem_14_shr_mem_14_or_cse_pff;
  assign shr_mem_14_cns_dinb_shi0 = MUX_v_64_2_2(dout_14_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_14_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_14_and_3_cse_pff);
  assign shr_mem_14_cns_addra_shi1 = shr_mem_14_shr_mem_14_mux_2_cse_pff;
  assign shr_mem_14_and_5_cse_pff = shr_mem_14_cns_S1_pff & shr_mem_14_xor_1_rmff;
  assign shr_mem_14_shr_mem_14_mux_2_cse_pff = MUX_v_8_2_2(dout_14_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_14_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_14_and_5_cse_pff);
  assign shr_mem_14_cns_addrb_shi1 = shr_mem_14_shr_mem_14_mux_2_cse_pff;
  assign shr_mem_14_cns_csa_n_shi1 = shr_mem_14_shr_mem_14_or_1_cse_pff;
  assign shr_mem_14_mux_7_nl = MUX_s_1_2_2(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_14_and_5_cse_pff);
  assign shr_mem_14_shr_mem_14_or_1_cse_pff = (shr_mem_14_mux_7_nl) | (~((shr_mem_14_cns_S0_pff
      & shr_mem_14_xor_rmff) | shr_mem_14_and_5_cse_pff));
  assign shr_mem_14_cns_csb_n_shi1 = shr_mem_14_shr_mem_14_or_1_cse_pff;
  assign shr_mem_14_cns_dinb_shi1 = MUX_v_64_2_2(dout_14_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_14_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_14_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_14_cns_ppidx <= 1'b0;
      shr_mem_14_cns_ppown <= 2'b0;
      shr_mem_14_cns_ppidx_1 <= 1'b0;
      shr_mem_14_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_14_cns_ppidx <= shr_mem_14_xor_rmff;
      shr_mem_14_cns_ppown <= shr_mem_14_acc_rmff;
      shr_mem_14_cns_ppidx_1 <= shr_mem_14_xor_1_rmff;
      shr_mem_14_cns_ppown_1 <= shr_mem_14_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffefnCNP13_cns_bctl
// ------------------------------------------------------------------


module double_buffefnCNP13_cns_bctl (
  clk, rst, dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_13_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_13_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_13_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_13_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_13_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_13_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_13_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_13_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_13_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_13_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_13_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_13_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_13_cns_S0, shr_mem_13_cns_R0, shr_mem_13_cns_S1, shr_mem_13_cns_R1,
      shr_mem_13_cns_addra_shi0, shr_mem_13_cns_addra_shi1, shr_mem_13_cns_addrb_shi0,
      shr_mem_13_cns_addrb_shi1, shr_mem_13_cns_csa_n_shi0, shr_mem_13_cns_csa_n_shi1,
      shr_mem_13_cns_csb_n_shi0, shr_mem_13_cns_csb_n_shi1, shr_mem_13_cns_dinb_shi0,
      shr_mem_13_cns_dinb_shi1, shr_mem_13_cns_douta_sho0, shr_mem_13_cns_douta_sho1,
      shr_mem_13_cns_S1_pff, din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_13_cns_S0_pff
);
  input clk;
  input rst;
  input dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_13_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_13_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_13_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_13_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_13_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_13_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_13_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_13_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_13_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_13_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_13_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_13_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_13_cns_S0;
  input shr_mem_13_cns_R0;
  output shr_mem_13_cns_S1;
  input shr_mem_13_cns_R1;
  output [7:0] shr_mem_13_cns_addra_shi0;
  output [7:0] shr_mem_13_cns_addra_shi1;
  output [7:0] shr_mem_13_cns_addrb_shi0;
  output [7:0] shr_mem_13_cns_addrb_shi1;
  output shr_mem_13_cns_csa_n_shi0;
  output shr_mem_13_cns_csa_n_shi1;
  output shr_mem_13_cns_csb_n_shi0;
  output shr_mem_13_cns_csb_n_shi1;
  output [63:0] shr_mem_13_cns_dinb_shi0;
  output [63:0] shr_mem_13_cns_dinb_shi1;
  input [63:0] shr_mem_13_cns_douta_sho0;
  input [63:0] shr_mem_13_cns_douta_sho1;
  output shr_mem_13_cns_S1_pff;
  input din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_13_cns_S0_pff;


  // Interconnect Declarations
  reg dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_13_cns_PC0;
  reg shr_mem_13_cns_ppidx;
  reg [1:0] shr_mem_13_cns_ppown;
  wire shr_mem_13_cns_PC1;
  reg shr_mem_13_cns_ppidx_1;
  reg [1:0] shr_mem_13_cns_ppown_1;
  wire [7:0] shr_mem_13_shr_mem_13_mux_3_cse_pff;
  wire shr_mem_13_and_3_cse_pff;
  wire [1:0] shr_mem_13_acc_1_rmff;
  wire [3:0] nl_shr_mem_13_acc_1_rmff;
  wire shr_mem_13_xor_1_rmff;
  wire shr_mem_13_shr_mem_13_or_cse_pff;
  wire [1:0] shr_mem_13_acc_rmff;
  wire [3:0] nl_shr_mem_13_acc_rmff;
  wire shr_mem_13_xor_rmff;
  wire [7:0] shr_mem_13_shr_mem_13_mux_2_cse_pff;
  wire shr_mem_13_and_5_cse_pff;
  wire shr_mem_13_shr_mem_13_or_1_cse_pff;

  wire[0:0] shr_mem_13_mux_6_nl;
  wire[0:0] shr_mem_13_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_13_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_13_cns_R0;
  assign din_13_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_13_cns_R1;
  assign shr_mem_13_xor_rmff = shr_mem_13_cns_ppidx ^ shr_mem_13_cns_PC0;
  assign nl_shr_mem_13_acc_rmff = shr_mem_13_cns_ppown + conv_u2u_1_2(shr_mem_13_cns_PC0)
      + conv_s2u_1_2(shr_mem_13_cns_PC1);
  assign shr_mem_13_acc_rmff = nl_shr_mem_13_acc_rmff[1:0];
  assign shr_mem_13_cns_PC0 = shr_mem_13_cns_S0 & dout_13_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_13_xor_1_rmff = shr_mem_13_cns_ppidx_1 ^ shr_mem_13_cns_PC1;
  assign nl_shr_mem_13_acc_1_rmff = shr_mem_13_cns_ppown_1 + conv_u2u_1_2(shr_mem_13_cns_PC1)
      + conv_s2u_1_2(shr_mem_13_cns_PC0);
  assign shr_mem_13_acc_1_rmff = nl_shr_mem_13_acc_1_rmff[1:0];
  assign shr_mem_13_cns_PC1 = shr_mem_13_cns_S1 & din_13_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_13_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_13_cns_douta_sho0,
      shr_mem_13_cns_douta_sho1, shr_mem_13_cns_ppidx);
  assign din_13_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_13_cns_douta_sho0,
      shr_mem_13_cns_douta_sho1, shr_mem_13_cns_ppidx_1);
  assign shr_mem_13_cns_addra_shi0 = shr_mem_13_shr_mem_13_mux_3_cse_pff;
  assign shr_mem_13_cns_S1 = (shr_mem_13_cns_ppown_1!=2'b00);
  assign shr_mem_13_cns_S1_pff = (shr_mem_13_acc_1_rmff!=2'b00);
  assign shr_mem_13_and_3_cse_pff = shr_mem_13_cns_S1_pff & (~ shr_mem_13_xor_1_rmff);
  assign shr_mem_13_shr_mem_13_mux_3_cse_pff = MUX_v_8_2_2(dout_13_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_13_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_13_and_3_cse_pff);
  assign shr_mem_13_cns_addrb_shi0 = shr_mem_13_shr_mem_13_mux_3_cse_pff;
  assign shr_mem_13_cns_csa_n_shi0 = shr_mem_13_shr_mem_13_or_cse_pff;
  assign din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_13_cns_S0 = ~((shr_mem_13_cns_ppown==2'b10));
  assign shr_mem_13_cns_S0_pff = ~((shr_mem_13_acc_rmff==2'b10));
  assign shr_mem_13_mux_6_nl = MUX_s_1_2_2(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_13_and_3_cse_pff);
  assign shr_mem_13_shr_mem_13_or_cse_pff = (shr_mem_13_mux_6_nl) | (~((shr_mem_13_cns_S0_pff
      & (~ shr_mem_13_xor_rmff)) | shr_mem_13_and_3_cse_pff));
  assign shr_mem_13_cns_csb_n_shi0 = shr_mem_13_shr_mem_13_or_cse_pff;
  assign shr_mem_13_cns_dinb_shi0 = MUX_v_64_2_2(dout_13_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_13_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_13_and_3_cse_pff);
  assign shr_mem_13_cns_addra_shi1 = shr_mem_13_shr_mem_13_mux_2_cse_pff;
  assign shr_mem_13_and_5_cse_pff = shr_mem_13_cns_S1_pff & shr_mem_13_xor_1_rmff;
  assign shr_mem_13_shr_mem_13_mux_2_cse_pff = MUX_v_8_2_2(dout_13_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_13_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_13_and_5_cse_pff);
  assign shr_mem_13_cns_addrb_shi1 = shr_mem_13_shr_mem_13_mux_2_cse_pff;
  assign shr_mem_13_cns_csa_n_shi1 = shr_mem_13_shr_mem_13_or_1_cse_pff;
  assign shr_mem_13_mux_7_nl = MUX_s_1_2_2(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_13_and_5_cse_pff);
  assign shr_mem_13_shr_mem_13_or_1_cse_pff = (shr_mem_13_mux_7_nl) | (~((shr_mem_13_cns_S0_pff
      & shr_mem_13_xor_rmff) | shr_mem_13_and_5_cse_pff));
  assign shr_mem_13_cns_csb_n_shi1 = shr_mem_13_shr_mem_13_or_1_cse_pff;
  assign shr_mem_13_cns_dinb_shi1 = MUX_v_64_2_2(dout_13_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_13_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_13_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_13_cns_ppidx <= 1'b0;
      shr_mem_13_cns_ppown <= 2'b0;
      shr_mem_13_cns_ppidx_1 <= 1'b0;
      shr_mem_13_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_13_cns_ppidx <= shr_mem_13_xor_rmff;
      shr_mem_13_cns_ppown <= shr_mem_13_acc_rmff;
      shr_mem_13_cns_ppidx_1 <= shr_mem_13_xor_1_rmff;
      shr_mem_13_cns_ppown_1 <= shr_mem_13_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffefnCNP12_cns_bctl
// ------------------------------------------------------------------


module double_buffefnCNP12_cns_bctl (
  clk, rst, dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_12_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_12_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_12_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_12_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_12_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_12_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_12_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_12_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_12_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_12_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_12_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_12_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_12_cns_S0, shr_mem_12_cns_R0, shr_mem_12_cns_S1, shr_mem_12_cns_R1,
      shr_mem_12_cns_addra_shi0, shr_mem_12_cns_addra_shi1, shr_mem_12_cns_addrb_shi0,
      shr_mem_12_cns_addrb_shi1, shr_mem_12_cns_csa_n_shi0, shr_mem_12_cns_csa_n_shi1,
      shr_mem_12_cns_csb_n_shi0, shr_mem_12_cns_csb_n_shi1, shr_mem_12_cns_dinb_shi0,
      shr_mem_12_cns_dinb_shi1, shr_mem_12_cns_douta_sho0, shr_mem_12_cns_douta_sho1,
      shr_mem_12_cns_S1_pff, din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_12_cns_S0_pff
);
  input clk;
  input rst;
  input dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_12_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_12_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_12_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_12_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_12_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_12_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_12_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_12_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_12_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_12_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_12_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_12_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_12_cns_S0;
  input shr_mem_12_cns_R0;
  output shr_mem_12_cns_S1;
  input shr_mem_12_cns_R1;
  output [7:0] shr_mem_12_cns_addra_shi0;
  output [7:0] shr_mem_12_cns_addra_shi1;
  output [7:0] shr_mem_12_cns_addrb_shi0;
  output [7:0] shr_mem_12_cns_addrb_shi1;
  output shr_mem_12_cns_csa_n_shi0;
  output shr_mem_12_cns_csa_n_shi1;
  output shr_mem_12_cns_csb_n_shi0;
  output shr_mem_12_cns_csb_n_shi1;
  output [63:0] shr_mem_12_cns_dinb_shi0;
  output [63:0] shr_mem_12_cns_dinb_shi1;
  input [63:0] shr_mem_12_cns_douta_sho0;
  input [63:0] shr_mem_12_cns_douta_sho1;
  output shr_mem_12_cns_S1_pff;
  input din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_12_cns_S0_pff;


  // Interconnect Declarations
  reg dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_12_cns_PC0;
  reg shr_mem_12_cns_ppidx;
  reg [1:0] shr_mem_12_cns_ppown;
  wire shr_mem_12_cns_PC1;
  reg shr_mem_12_cns_ppidx_1;
  reg [1:0] shr_mem_12_cns_ppown_1;
  wire [7:0] shr_mem_12_shr_mem_12_mux_3_cse_pff;
  wire shr_mem_12_and_3_cse_pff;
  wire [1:0] shr_mem_12_acc_1_rmff;
  wire [3:0] nl_shr_mem_12_acc_1_rmff;
  wire shr_mem_12_xor_1_rmff;
  wire shr_mem_12_shr_mem_12_or_cse_pff;
  wire [1:0] shr_mem_12_acc_rmff;
  wire [3:0] nl_shr_mem_12_acc_rmff;
  wire shr_mem_12_xor_rmff;
  wire [7:0] shr_mem_12_shr_mem_12_mux_2_cse_pff;
  wire shr_mem_12_and_5_cse_pff;
  wire shr_mem_12_shr_mem_12_or_1_cse_pff;

  wire[0:0] shr_mem_12_mux_6_nl;
  wire[0:0] shr_mem_12_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_12_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_12_cns_R0;
  assign din_12_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_12_cns_R1;
  assign shr_mem_12_xor_rmff = shr_mem_12_cns_ppidx ^ shr_mem_12_cns_PC0;
  assign nl_shr_mem_12_acc_rmff = shr_mem_12_cns_ppown + conv_u2u_1_2(shr_mem_12_cns_PC0)
      + conv_s2u_1_2(shr_mem_12_cns_PC1);
  assign shr_mem_12_acc_rmff = nl_shr_mem_12_acc_rmff[1:0];
  assign shr_mem_12_cns_PC0 = shr_mem_12_cns_S0 & dout_12_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_12_xor_1_rmff = shr_mem_12_cns_ppidx_1 ^ shr_mem_12_cns_PC1;
  assign nl_shr_mem_12_acc_1_rmff = shr_mem_12_cns_ppown_1 + conv_u2u_1_2(shr_mem_12_cns_PC1)
      + conv_s2u_1_2(shr_mem_12_cns_PC0);
  assign shr_mem_12_acc_1_rmff = nl_shr_mem_12_acc_1_rmff[1:0];
  assign shr_mem_12_cns_PC1 = shr_mem_12_cns_S1 & din_12_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_12_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_12_cns_douta_sho0,
      shr_mem_12_cns_douta_sho1, shr_mem_12_cns_ppidx);
  assign din_12_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_12_cns_douta_sho0,
      shr_mem_12_cns_douta_sho1, shr_mem_12_cns_ppidx_1);
  assign shr_mem_12_cns_addra_shi0 = shr_mem_12_shr_mem_12_mux_3_cse_pff;
  assign shr_mem_12_cns_S1 = (shr_mem_12_cns_ppown_1!=2'b00);
  assign shr_mem_12_cns_S1_pff = (shr_mem_12_acc_1_rmff!=2'b00);
  assign shr_mem_12_and_3_cse_pff = shr_mem_12_cns_S1_pff & (~ shr_mem_12_xor_1_rmff);
  assign shr_mem_12_shr_mem_12_mux_3_cse_pff = MUX_v_8_2_2(dout_12_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_12_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_12_and_3_cse_pff);
  assign shr_mem_12_cns_addrb_shi0 = shr_mem_12_shr_mem_12_mux_3_cse_pff;
  assign shr_mem_12_cns_csa_n_shi0 = shr_mem_12_shr_mem_12_or_cse_pff;
  assign din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_12_cns_S0 = ~((shr_mem_12_cns_ppown==2'b10));
  assign shr_mem_12_cns_S0_pff = ~((shr_mem_12_acc_rmff==2'b10));
  assign shr_mem_12_mux_6_nl = MUX_s_1_2_2(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_12_and_3_cse_pff);
  assign shr_mem_12_shr_mem_12_or_cse_pff = (shr_mem_12_mux_6_nl) | (~((shr_mem_12_cns_S0_pff
      & (~ shr_mem_12_xor_rmff)) | shr_mem_12_and_3_cse_pff));
  assign shr_mem_12_cns_csb_n_shi0 = shr_mem_12_shr_mem_12_or_cse_pff;
  assign shr_mem_12_cns_dinb_shi0 = MUX_v_64_2_2(dout_12_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_12_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_12_and_3_cse_pff);
  assign shr_mem_12_cns_addra_shi1 = shr_mem_12_shr_mem_12_mux_2_cse_pff;
  assign shr_mem_12_and_5_cse_pff = shr_mem_12_cns_S1_pff & shr_mem_12_xor_1_rmff;
  assign shr_mem_12_shr_mem_12_mux_2_cse_pff = MUX_v_8_2_2(dout_12_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_12_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_12_and_5_cse_pff);
  assign shr_mem_12_cns_addrb_shi1 = shr_mem_12_shr_mem_12_mux_2_cse_pff;
  assign shr_mem_12_cns_csa_n_shi1 = shr_mem_12_shr_mem_12_or_1_cse_pff;
  assign shr_mem_12_mux_7_nl = MUX_s_1_2_2(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_12_and_5_cse_pff);
  assign shr_mem_12_shr_mem_12_or_1_cse_pff = (shr_mem_12_mux_7_nl) | (~((shr_mem_12_cns_S0_pff
      & shr_mem_12_xor_rmff) | shr_mem_12_and_5_cse_pff));
  assign shr_mem_12_cns_csb_n_shi1 = shr_mem_12_shr_mem_12_or_1_cse_pff;
  assign shr_mem_12_cns_dinb_shi1 = MUX_v_64_2_2(dout_12_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_12_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_12_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_12_cns_ppidx <= 1'b0;
      shr_mem_12_cns_ppown <= 2'b0;
      shr_mem_12_cns_ppidx_1 <= 1'b0;
      shr_mem_12_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_12_cns_ppidx <= shr_mem_12_xor_rmff;
      shr_mem_12_cns_ppown <= shr_mem_12_acc_rmff;
      shr_mem_12_cns_ppidx_1 <= shr_mem_12_xor_1_rmff;
      shr_mem_12_cns_ppown_1 <= shr_mem_12_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffefnCNP11_cns_bctl
// ------------------------------------------------------------------


module double_buffefnCNP11_cns_bctl (
  clk, rst, dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_11_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_11_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_11_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_11_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_11_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_11_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_11_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_11_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_11_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_11_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_11_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_11_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_11_cns_S0, shr_mem_11_cns_R0, shr_mem_11_cns_S1, shr_mem_11_cns_R1,
      shr_mem_11_cns_addra_shi0, shr_mem_11_cns_addra_shi1, shr_mem_11_cns_addrb_shi0,
      shr_mem_11_cns_addrb_shi1, shr_mem_11_cns_csa_n_shi0, shr_mem_11_cns_csa_n_shi1,
      shr_mem_11_cns_csb_n_shi0, shr_mem_11_cns_csb_n_shi1, shr_mem_11_cns_dinb_shi0,
      shr_mem_11_cns_dinb_shi1, shr_mem_11_cns_douta_sho0, shr_mem_11_cns_douta_sho1,
      shr_mem_11_cns_S1_pff, din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_11_cns_S0_pff
);
  input clk;
  input rst;
  input dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_11_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_11_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_11_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_11_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_11_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_11_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_11_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_11_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_11_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_11_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_11_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_11_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_11_cns_S0;
  input shr_mem_11_cns_R0;
  output shr_mem_11_cns_S1;
  input shr_mem_11_cns_R1;
  output [7:0] shr_mem_11_cns_addra_shi0;
  output [7:0] shr_mem_11_cns_addra_shi1;
  output [7:0] shr_mem_11_cns_addrb_shi0;
  output [7:0] shr_mem_11_cns_addrb_shi1;
  output shr_mem_11_cns_csa_n_shi0;
  output shr_mem_11_cns_csa_n_shi1;
  output shr_mem_11_cns_csb_n_shi0;
  output shr_mem_11_cns_csb_n_shi1;
  output [63:0] shr_mem_11_cns_dinb_shi0;
  output [63:0] shr_mem_11_cns_dinb_shi1;
  input [63:0] shr_mem_11_cns_douta_sho0;
  input [63:0] shr_mem_11_cns_douta_sho1;
  output shr_mem_11_cns_S1_pff;
  input din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_11_cns_S0_pff;


  // Interconnect Declarations
  reg dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_11_cns_PC0;
  reg shr_mem_11_cns_ppidx;
  reg [1:0] shr_mem_11_cns_ppown;
  wire shr_mem_11_cns_PC1;
  reg shr_mem_11_cns_ppidx_1;
  reg [1:0] shr_mem_11_cns_ppown_1;
  wire [7:0] shr_mem_11_shr_mem_11_mux_3_cse_pff;
  wire shr_mem_11_and_3_cse_pff;
  wire [1:0] shr_mem_11_acc_1_rmff;
  wire [3:0] nl_shr_mem_11_acc_1_rmff;
  wire shr_mem_11_xor_1_rmff;
  wire shr_mem_11_shr_mem_11_or_cse_pff;
  wire [1:0] shr_mem_11_acc_rmff;
  wire [3:0] nl_shr_mem_11_acc_rmff;
  wire shr_mem_11_xor_rmff;
  wire [7:0] shr_mem_11_shr_mem_11_mux_2_cse_pff;
  wire shr_mem_11_and_5_cse_pff;
  wire shr_mem_11_shr_mem_11_or_1_cse_pff;

  wire[0:0] shr_mem_11_mux_6_nl;
  wire[0:0] shr_mem_11_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_11_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_11_cns_R0;
  assign din_11_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_11_cns_R1;
  assign shr_mem_11_xor_rmff = shr_mem_11_cns_ppidx ^ shr_mem_11_cns_PC0;
  assign nl_shr_mem_11_acc_rmff = shr_mem_11_cns_ppown + conv_u2u_1_2(shr_mem_11_cns_PC0)
      + conv_s2u_1_2(shr_mem_11_cns_PC1);
  assign shr_mem_11_acc_rmff = nl_shr_mem_11_acc_rmff[1:0];
  assign shr_mem_11_cns_PC0 = shr_mem_11_cns_S0 & dout_11_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_11_xor_1_rmff = shr_mem_11_cns_ppidx_1 ^ shr_mem_11_cns_PC1;
  assign nl_shr_mem_11_acc_1_rmff = shr_mem_11_cns_ppown_1 + conv_u2u_1_2(shr_mem_11_cns_PC1)
      + conv_s2u_1_2(shr_mem_11_cns_PC0);
  assign shr_mem_11_acc_1_rmff = nl_shr_mem_11_acc_1_rmff[1:0];
  assign shr_mem_11_cns_PC1 = shr_mem_11_cns_S1 & din_11_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_11_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_11_cns_douta_sho0,
      shr_mem_11_cns_douta_sho1, shr_mem_11_cns_ppidx);
  assign din_11_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_11_cns_douta_sho0,
      shr_mem_11_cns_douta_sho1, shr_mem_11_cns_ppidx_1);
  assign shr_mem_11_cns_addra_shi0 = shr_mem_11_shr_mem_11_mux_3_cse_pff;
  assign shr_mem_11_cns_S1 = (shr_mem_11_cns_ppown_1!=2'b00);
  assign shr_mem_11_cns_S1_pff = (shr_mem_11_acc_1_rmff!=2'b00);
  assign shr_mem_11_and_3_cse_pff = shr_mem_11_cns_S1_pff & (~ shr_mem_11_xor_1_rmff);
  assign shr_mem_11_shr_mem_11_mux_3_cse_pff = MUX_v_8_2_2(dout_11_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_11_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_11_and_3_cse_pff);
  assign shr_mem_11_cns_addrb_shi0 = shr_mem_11_shr_mem_11_mux_3_cse_pff;
  assign shr_mem_11_cns_csa_n_shi0 = shr_mem_11_shr_mem_11_or_cse_pff;
  assign din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_11_cns_S0 = ~((shr_mem_11_cns_ppown==2'b10));
  assign shr_mem_11_cns_S0_pff = ~((shr_mem_11_acc_rmff==2'b10));
  assign shr_mem_11_mux_6_nl = MUX_s_1_2_2(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_11_and_3_cse_pff);
  assign shr_mem_11_shr_mem_11_or_cse_pff = (shr_mem_11_mux_6_nl) | (~((shr_mem_11_cns_S0_pff
      & (~ shr_mem_11_xor_rmff)) | shr_mem_11_and_3_cse_pff));
  assign shr_mem_11_cns_csb_n_shi0 = shr_mem_11_shr_mem_11_or_cse_pff;
  assign shr_mem_11_cns_dinb_shi0 = MUX_v_64_2_2(dout_11_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_11_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_11_and_3_cse_pff);
  assign shr_mem_11_cns_addra_shi1 = shr_mem_11_shr_mem_11_mux_2_cse_pff;
  assign shr_mem_11_and_5_cse_pff = shr_mem_11_cns_S1_pff & shr_mem_11_xor_1_rmff;
  assign shr_mem_11_shr_mem_11_mux_2_cse_pff = MUX_v_8_2_2(dout_11_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_11_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_11_and_5_cse_pff);
  assign shr_mem_11_cns_addrb_shi1 = shr_mem_11_shr_mem_11_mux_2_cse_pff;
  assign shr_mem_11_cns_csa_n_shi1 = shr_mem_11_shr_mem_11_or_1_cse_pff;
  assign shr_mem_11_mux_7_nl = MUX_s_1_2_2(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_11_and_5_cse_pff);
  assign shr_mem_11_shr_mem_11_or_1_cse_pff = (shr_mem_11_mux_7_nl) | (~((shr_mem_11_cns_S0_pff
      & shr_mem_11_xor_rmff) | shr_mem_11_and_5_cse_pff));
  assign shr_mem_11_cns_csb_n_shi1 = shr_mem_11_shr_mem_11_or_1_cse_pff;
  assign shr_mem_11_cns_dinb_shi1 = MUX_v_64_2_2(dout_11_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_11_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_11_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_11_cns_ppidx <= 1'b0;
      shr_mem_11_cns_ppown <= 2'b0;
      shr_mem_11_cns_ppidx_1 <= 1'b0;
      shr_mem_11_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_11_cns_ppidx <= shr_mem_11_xor_rmff;
      shr_mem_11_cns_ppown <= shr_mem_11_acc_rmff;
      shr_mem_11_cns_ppidx_1 <= shr_mem_11_xor_1_rmff;
      shr_mem_11_cns_ppown_1 <= shr_mem_11_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffefnCNP10_cns_bctl
// ------------------------------------------------------------------


module double_buffefnCNP10_cns_bctl (
  clk, rst, dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_10_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_10_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_10_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_10_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_10_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_10_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_10_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_10_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_10_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_10_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_10_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_10_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_10_cns_S0, shr_mem_10_cns_R0, shr_mem_10_cns_S1, shr_mem_10_cns_R1,
      shr_mem_10_cns_addra_shi0, shr_mem_10_cns_addra_shi1, shr_mem_10_cns_addrb_shi0,
      shr_mem_10_cns_addrb_shi1, shr_mem_10_cns_csa_n_shi0, shr_mem_10_cns_csa_n_shi1,
      shr_mem_10_cns_csb_n_shi0, shr_mem_10_cns_csb_n_shi1, shr_mem_10_cns_dinb_shi0,
      shr_mem_10_cns_dinb_shi1, shr_mem_10_cns_douta_sho0, shr_mem_10_cns_douta_sho1,
      shr_mem_10_cns_S1_pff, din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_10_cns_S0_pff
);
  input clk;
  input rst;
  input dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_10_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_10_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_10_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_10_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_10_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_10_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_10_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_10_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_10_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_10_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_10_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_10_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_10_cns_S0;
  input shr_mem_10_cns_R0;
  output shr_mem_10_cns_S1;
  input shr_mem_10_cns_R1;
  output [7:0] shr_mem_10_cns_addra_shi0;
  output [7:0] shr_mem_10_cns_addra_shi1;
  output [7:0] shr_mem_10_cns_addrb_shi0;
  output [7:0] shr_mem_10_cns_addrb_shi1;
  output shr_mem_10_cns_csa_n_shi0;
  output shr_mem_10_cns_csa_n_shi1;
  output shr_mem_10_cns_csb_n_shi0;
  output shr_mem_10_cns_csb_n_shi1;
  output [63:0] shr_mem_10_cns_dinb_shi0;
  output [63:0] shr_mem_10_cns_dinb_shi1;
  input [63:0] shr_mem_10_cns_douta_sho0;
  input [63:0] shr_mem_10_cns_douta_sho1;
  output shr_mem_10_cns_S1_pff;
  input din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_10_cns_S0_pff;


  // Interconnect Declarations
  reg dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_10_cns_PC0;
  reg shr_mem_10_cns_ppidx;
  reg [1:0] shr_mem_10_cns_ppown;
  wire shr_mem_10_cns_PC1;
  reg shr_mem_10_cns_ppidx_1;
  reg [1:0] shr_mem_10_cns_ppown_1;
  wire [7:0] shr_mem_10_shr_mem_10_mux_3_cse_pff;
  wire shr_mem_10_and_3_cse_pff;
  wire [1:0] shr_mem_10_acc_1_rmff;
  wire [3:0] nl_shr_mem_10_acc_1_rmff;
  wire shr_mem_10_xor_1_rmff;
  wire shr_mem_10_shr_mem_10_or_cse_pff;
  wire [1:0] shr_mem_10_acc_rmff;
  wire [3:0] nl_shr_mem_10_acc_rmff;
  wire shr_mem_10_xor_rmff;
  wire [7:0] shr_mem_10_shr_mem_10_mux_2_cse_pff;
  wire shr_mem_10_and_5_cse_pff;
  wire shr_mem_10_shr_mem_10_or_1_cse_pff;

  wire[0:0] shr_mem_10_mux_6_nl;
  wire[0:0] shr_mem_10_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_10_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_10_cns_R0;
  assign din_10_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_10_cns_R1;
  assign shr_mem_10_xor_rmff = shr_mem_10_cns_ppidx ^ shr_mem_10_cns_PC0;
  assign nl_shr_mem_10_acc_rmff = shr_mem_10_cns_ppown + conv_u2u_1_2(shr_mem_10_cns_PC0)
      + conv_s2u_1_2(shr_mem_10_cns_PC1);
  assign shr_mem_10_acc_rmff = nl_shr_mem_10_acc_rmff[1:0];
  assign shr_mem_10_cns_PC0 = shr_mem_10_cns_S0 & dout_10_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_10_xor_1_rmff = shr_mem_10_cns_ppidx_1 ^ shr_mem_10_cns_PC1;
  assign nl_shr_mem_10_acc_1_rmff = shr_mem_10_cns_ppown_1 + conv_u2u_1_2(shr_mem_10_cns_PC1)
      + conv_s2u_1_2(shr_mem_10_cns_PC0);
  assign shr_mem_10_acc_1_rmff = nl_shr_mem_10_acc_1_rmff[1:0];
  assign shr_mem_10_cns_PC1 = shr_mem_10_cns_S1 & din_10_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_10_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_10_cns_douta_sho0,
      shr_mem_10_cns_douta_sho1, shr_mem_10_cns_ppidx);
  assign din_10_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_10_cns_douta_sho0,
      shr_mem_10_cns_douta_sho1, shr_mem_10_cns_ppidx_1);
  assign shr_mem_10_cns_addra_shi0 = shr_mem_10_shr_mem_10_mux_3_cse_pff;
  assign shr_mem_10_cns_S1 = (shr_mem_10_cns_ppown_1!=2'b00);
  assign shr_mem_10_cns_S1_pff = (shr_mem_10_acc_1_rmff!=2'b00);
  assign shr_mem_10_and_3_cse_pff = shr_mem_10_cns_S1_pff & (~ shr_mem_10_xor_1_rmff);
  assign shr_mem_10_shr_mem_10_mux_3_cse_pff = MUX_v_8_2_2(dout_10_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_10_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_10_and_3_cse_pff);
  assign shr_mem_10_cns_addrb_shi0 = shr_mem_10_shr_mem_10_mux_3_cse_pff;
  assign shr_mem_10_cns_csa_n_shi0 = shr_mem_10_shr_mem_10_or_cse_pff;
  assign din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_10_cns_S0 = ~((shr_mem_10_cns_ppown==2'b10));
  assign shr_mem_10_cns_S0_pff = ~((shr_mem_10_acc_rmff==2'b10));
  assign shr_mem_10_mux_6_nl = MUX_s_1_2_2(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_10_and_3_cse_pff);
  assign shr_mem_10_shr_mem_10_or_cse_pff = (shr_mem_10_mux_6_nl) | (~((shr_mem_10_cns_S0_pff
      & (~ shr_mem_10_xor_rmff)) | shr_mem_10_and_3_cse_pff));
  assign shr_mem_10_cns_csb_n_shi0 = shr_mem_10_shr_mem_10_or_cse_pff;
  assign shr_mem_10_cns_dinb_shi0 = MUX_v_64_2_2(dout_10_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_10_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_10_and_3_cse_pff);
  assign shr_mem_10_cns_addra_shi1 = shr_mem_10_shr_mem_10_mux_2_cse_pff;
  assign shr_mem_10_and_5_cse_pff = shr_mem_10_cns_S1_pff & shr_mem_10_xor_1_rmff;
  assign shr_mem_10_shr_mem_10_mux_2_cse_pff = MUX_v_8_2_2(dout_10_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_10_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_10_and_5_cse_pff);
  assign shr_mem_10_cns_addrb_shi1 = shr_mem_10_shr_mem_10_mux_2_cse_pff;
  assign shr_mem_10_cns_csa_n_shi1 = shr_mem_10_shr_mem_10_or_1_cse_pff;
  assign shr_mem_10_mux_7_nl = MUX_s_1_2_2(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_10_and_5_cse_pff);
  assign shr_mem_10_shr_mem_10_or_1_cse_pff = (shr_mem_10_mux_7_nl) | (~((shr_mem_10_cns_S0_pff
      & shr_mem_10_xor_rmff) | shr_mem_10_and_5_cse_pff));
  assign shr_mem_10_cns_csb_n_shi1 = shr_mem_10_shr_mem_10_or_1_cse_pff;
  assign shr_mem_10_cns_dinb_shi1 = MUX_v_64_2_2(dout_10_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_10_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_10_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_10_cns_ppidx <= 1'b0;
      shr_mem_10_cns_ppown <= 2'b0;
      shr_mem_10_cns_ppidx_1 <= 1'b0;
      shr_mem_10_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_10_cns_ppidx <= shr_mem_10_xor_rmff;
      shr_mem_10_cns_ppown <= shr_mem_10_acc_rmff;
      shr_mem_10_cns_ppidx_1 <= shr_mem_10_xor_1_rmff;
      shr_mem_10_cns_ppown_1 <= shr_mem_10_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeYeetf_9_cns_bctl
// ------------------------------------------------------------------


module double_buffeYeetf_9_cns_bctl (
  clk, rst, dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_9_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_9_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_9_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_9_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_9_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_9_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_9_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_9_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_9_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_9_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_9_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_9_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_9_cns_S0, shr_mem_9_cns_R0, shr_mem_9_cns_S1, shr_mem_9_cns_R1, shr_mem_9_cns_addra_shi0,
      shr_mem_9_cns_addra_shi1, shr_mem_9_cns_addrb_shi0, shr_mem_9_cns_addrb_shi1,
      shr_mem_9_cns_csa_n_shi0, shr_mem_9_cns_csa_n_shi1, shr_mem_9_cns_csb_n_shi0,
      shr_mem_9_cns_csb_n_shi1, shr_mem_9_cns_dinb_shi0, shr_mem_9_cns_dinb_shi1,
      shr_mem_9_cns_douta_sho0, shr_mem_9_cns_douta_sho1, shr_mem_9_cns_S1_pff, din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_9_cns_S0_pff
);
  input clk;
  input rst;
  input dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_9_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_9_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_9_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_9_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_9_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_9_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_9_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_9_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_9_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_9_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_9_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_9_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_9_cns_S0;
  input shr_mem_9_cns_R0;
  output shr_mem_9_cns_S1;
  input shr_mem_9_cns_R1;
  output [7:0] shr_mem_9_cns_addra_shi0;
  output [7:0] shr_mem_9_cns_addra_shi1;
  output [7:0] shr_mem_9_cns_addrb_shi0;
  output [7:0] shr_mem_9_cns_addrb_shi1;
  output shr_mem_9_cns_csa_n_shi0;
  output shr_mem_9_cns_csa_n_shi1;
  output shr_mem_9_cns_csb_n_shi0;
  output shr_mem_9_cns_csb_n_shi1;
  output [63:0] shr_mem_9_cns_dinb_shi0;
  output [63:0] shr_mem_9_cns_dinb_shi1;
  input [63:0] shr_mem_9_cns_douta_sho0;
  input [63:0] shr_mem_9_cns_douta_sho1;
  output shr_mem_9_cns_S1_pff;
  input din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_9_cns_S0_pff;


  // Interconnect Declarations
  reg dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_9_cns_PC0;
  reg shr_mem_9_cns_ppidx;
  reg [1:0] shr_mem_9_cns_ppown;
  wire shr_mem_9_cns_PC1;
  reg shr_mem_9_cns_ppidx_1;
  reg [1:0] shr_mem_9_cns_ppown_1;
  wire [7:0] shr_mem_9_shr_mem_9_mux_3_cse_pff;
  wire shr_mem_9_and_3_cse_pff;
  wire [1:0] shr_mem_9_acc_1_rmff;
  wire [3:0] nl_shr_mem_9_acc_1_rmff;
  wire shr_mem_9_xor_1_rmff;
  wire shr_mem_9_shr_mem_9_or_cse_pff;
  wire [1:0] shr_mem_9_acc_rmff;
  wire [3:0] nl_shr_mem_9_acc_rmff;
  wire shr_mem_9_xor_rmff;
  wire [7:0] shr_mem_9_shr_mem_9_mux_2_cse_pff;
  wire shr_mem_9_and_5_cse_pff;
  wire shr_mem_9_shr_mem_9_or_1_cse_pff;

  wire[0:0] shr_mem_9_mux_6_nl;
  wire[0:0] shr_mem_9_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_9_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_9_cns_R0;
  assign din_9_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_9_cns_R1;
  assign shr_mem_9_xor_rmff = shr_mem_9_cns_ppidx ^ shr_mem_9_cns_PC0;
  assign nl_shr_mem_9_acc_rmff = shr_mem_9_cns_ppown + conv_u2u_1_2(shr_mem_9_cns_PC0)
      + conv_s2u_1_2(shr_mem_9_cns_PC1);
  assign shr_mem_9_acc_rmff = nl_shr_mem_9_acc_rmff[1:0];
  assign shr_mem_9_cns_PC0 = shr_mem_9_cns_S0 & dout_9_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_9_xor_1_rmff = shr_mem_9_cns_ppidx_1 ^ shr_mem_9_cns_PC1;
  assign nl_shr_mem_9_acc_1_rmff = shr_mem_9_cns_ppown_1 + conv_u2u_1_2(shr_mem_9_cns_PC1)
      + conv_s2u_1_2(shr_mem_9_cns_PC0);
  assign shr_mem_9_acc_1_rmff = nl_shr_mem_9_acc_1_rmff[1:0];
  assign shr_mem_9_cns_PC1 = shr_mem_9_cns_S1 & din_9_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_9_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_9_cns_douta_sho0,
      shr_mem_9_cns_douta_sho1, shr_mem_9_cns_ppidx);
  assign din_9_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_9_cns_douta_sho0,
      shr_mem_9_cns_douta_sho1, shr_mem_9_cns_ppidx_1);
  assign shr_mem_9_cns_addra_shi0 = shr_mem_9_shr_mem_9_mux_3_cse_pff;
  assign shr_mem_9_cns_S1 = (shr_mem_9_cns_ppown_1!=2'b00);
  assign shr_mem_9_cns_S1_pff = (shr_mem_9_acc_1_rmff!=2'b00);
  assign shr_mem_9_and_3_cse_pff = shr_mem_9_cns_S1_pff & (~ shr_mem_9_xor_1_rmff);
  assign shr_mem_9_shr_mem_9_mux_3_cse_pff = MUX_v_8_2_2(dout_9_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_9_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_9_and_3_cse_pff);
  assign shr_mem_9_cns_addrb_shi0 = shr_mem_9_shr_mem_9_mux_3_cse_pff;
  assign shr_mem_9_cns_csa_n_shi0 = shr_mem_9_shr_mem_9_or_cse_pff;
  assign din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_9_cns_S0 = ~((shr_mem_9_cns_ppown==2'b10));
  assign shr_mem_9_cns_S0_pff = ~((shr_mem_9_acc_rmff==2'b10));
  assign shr_mem_9_mux_6_nl = MUX_s_1_2_2(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_9_and_3_cse_pff);
  assign shr_mem_9_shr_mem_9_or_cse_pff = (shr_mem_9_mux_6_nl) | (~((shr_mem_9_cns_S0_pff
      & (~ shr_mem_9_xor_rmff)) | shr_mem_9_and_3_cse_pff));
  assign shr_mem_9_cns_csb_n_shi0 = shr_mem_9_shr_mem_9_or_cse_pff;
  assign shr_mem_9_cns_dinb_shi0 = MUX_v_64_2_2(dout_9_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_9_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_9_and_3_cse_pff);
  assign shr_mem_9_cns_addra_shi1 = shr_mem_9_shr_mem_9_mux_2_cse_pff;
  assign shr_mem_9_and_5_cse_pff = shr_mem_9_cns_S1_pff & shr_mem_9_xor_1_rmff;
  assign shr_mem_9_shr_mem_9_mux_2_cse_pff = MUX_v_8_2_2(dout_9_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_9_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_9_and_5_cse_pff);
  assign shr_mem_9_cns_addrb_shi1 = shr_mem_9_shr_mem_9_mux_2_cse_pff;
  assign shr_mem_9_cns_csa_n_shi1 = shr_mem_9_shr_mem_9_or_1_cse_pff;
  assign shr_mem_9_mux_7_nl = MUX_s_1_2_2(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_9_and_5_cse_pff);
  assign shr_mem_9_shr_mem_9_or_1_cse_pff = (shr_mem_9_mux_7_nl) | (~((shr_mem_9_cns_S0_pff
      & shr_mem_9_xor_rmff) | shr_mem_9_and_5_cse_pff));
  assign shr_mem_9_cns_csb_n_shi1 = shr_mem_9_shr_mem_9_or_1_cse_pff;
  assign shr_mem_9_cns_dinb_shi1 = MUX_v_64_2_2(dout_9_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_9_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_9_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_9_cns_ppidx <= 1'b0;
      shr_mem_9_cns_ppown <= 2'b0;
      shr_mem_9_cns_ppidx_1 <= 1'b0;
      shr_mem_9_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_9_cns_ppidx <= shr_mem_9_xor_rmff;
      shr_mem_9_cns_ppown <= shr_mem_9_acc_rmff;
      shr_mem_9_cns_ppidx_1 <= shr_mem_9_xor_1_rmff;
      shr_mem_9_cns_ppown_1 <= shr_mem_9_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeYeetf_8_cns_bctl
// ------------------------------------------------------------------


module double_buffeYeetf_8_cns_bctl (
  clk, rst, dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_8_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_8_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_8_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_8_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_8_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_8_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_8_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_8_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_8_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_8_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_8_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_8_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_8_cns_S0, shr_mem_8_cns_R0, shr_mem_8_cns_S1, shr_mem_8_cns_R1, shr_mem_8_cns_addra_shi0,
      shr_mem_8_cns_addra_shi1, shr_mem_8_cns_addrb_shi0, shr_mem_8_cns_addrb_shi1,
      shr_mem_8_cns_csa_n_shi0, shr_mem_8_cns_csa_n_shi1, shr_mem_8_cns_csb_n_shi0,
      shr_mem_8_cns_csb_n_shi1, shr_mem_8_cns_dinb_shi0, shr_mem_8_cns_dinb_shi1,
      shr_mem_8_cns_douta_sho0, shr_mem_8_cns_douta_sho1, shr_mem_8_cns_S1_pff, din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_8_cns_S0_pff
);
  input clk;
  input rst;
  input dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_8_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_8_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_8_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_8_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_8_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_8_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_8_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_8_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_8_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_8_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_8_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_8_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_8_cns_S0;
  input shr_mem_8_cns_R0;
  output shr_mem_8_cns_S1;
  input shr_mem_8_cns_R1;
  output [7:0] shr_mem_8_cns_addra_shi0;
  output [7:0] shr_mem_8_cns_addra_shi1;
  output [7:0] shr_mem_8_cns_addrb_shi0;
  output [7:0] shr_mem_8_cns_addrb_shi1;
  output shr_mem_8_cns_csa_n_shi0;
  output shr_mem_8_cns_csa_n_shi1;
  output shr_mem_8_cns_csb_n_shi0;
  output shr_mem_8_cns_csb_n_shi1;
  output [63:0] shr_mem_8_cns_dinb_shi0;
  output [63:0] shr_mem_8_cns_dinb_shi1;
  input [63:0] shr_mem_8_cns_douta_sho0;
  input [63:0] shr_mem_8_cns_douta_sho1;
  output shr_mem_8_cns_S1_pff;
  input din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_8_cns_S0_pff;


  // Interconnect Declarations
  reg dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_8_cns_PC0;
  reg shr_mem_8_cns_ppidx;
  reg [1:0] shr_mem_8_cns_ppown;
  wire shr_mem_8_cns_PC1;
  reg shr_mem_8_cns_ppidx_1;
  reg [1:0] shr_mem_8_cns_ppown_1;
  wire [7:0] shr_mem_8_shr_mem_8_mux_3_cse_pff;
  wire shr_mem_8_and_3_cse_pff;
  wire [1:0] shr_mem_8_acc_1_rmff;
  wire [3:0] nl_shr_mem_8_acc_1_rmff;
  wire shr_mem_8_xor_1_rmff;
  wire shr_mem_8_shr_mem_8_or_cse_pff;
  wire [1:0] shr_mem_8_acc_rmff;
  wire [3:0] nl_shr_mem_8_acc_rmff;
  wire shr_mem_8_xor_rmff;
  wire [7:0] shr_mem_8_shr_mem_8_mux_2_cse_pff;
  wire shr_mem_8_and_5_cse_pff;
  wire shr_mem_8_shr_mem_8_or_1_cse_pff;

  wire[0:0] shr_mem_8_mux_6_nl;
  wire[0:0] shr_mem_8_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_8_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_8_cns_R0;
  assign din_8_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_8_cns_R1;
  assign shr_mem_8_xor_rmff = shr_mem_8_cns_ppidx ^ shr_mem_8_cns_PC0;
  assign nl_shr_mem_8_acc_rmff = shr_mem_8_cns_ppown + conv_u2u_1_2(shr_mem_8_cns_PC0)
      + conv_s2u_1_2(shr_mem_8_cns_PC1);
  assign shr_mem_8_acc_rmff = nl_shr_mem_8_acc_rmff[1:0];
  assign shr_mem_8_cns_PC0 = shr_mem_8_cns_S0 & dout_8_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_8_xor_1_rmff = shr_mem_8_cns_ppidx_1 ^ shr_mem_8_cns_PC1;
  assign nl_shr_mem_8_acc_1_rmff = shr_mem_8_cns_ppown_1 + conv_u2u_1_2(shr_mem_8_cns_PC1)
      + conv_s2u_1_2(shr_mem_8_cns_PC0);
  assign shr_mem_8_acc_1_rmff = nl_shr_mem_8_acc_1_rmff[1:0];
  assign shr_mem_8_cns_PC1 = shr_mem_8_cns_S1 & din_8_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_8_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_8_cns_douta_sho0,
      shr_mem_8_cns_douta_sho1, shr_mem_8_cns_ppidx);
  assign din_8_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_8_cns_douta_sho0,
      shr_mem_8_cns_douta_sho1, shr_mem_8_cns_ppidx_1);
  assign shr_mem_8_cns_addra_shi0 = shr_mem_8_shr_mem_8_mux_3_cse_pff;
  assign shr_mem_8_cns_S1 = (shr_mem_8_cns_ppown_1!=2'b00);
  assign shr_mem_8_cns_S1_pff = (shr_mem_8_acc_1_rmff!=2'b00);
  assign shr_mem_8_and_3_cse_pff = shr_mem_8_cns_S1_pff & (~ shr_mem_8_xor_1_rmff);
  assign shr_mem_8_shr_mem_8_mux_3_cse_pff = MUX_v_8_2_2(dout_8_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_8_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_8_and_3_cse_pff);
  assign shr_mem_8_cns_addrb_shi0 = shr_mem_8_shr_mem_8_mux_3_cse_pff;
  assign shr_mem_8_cns_csa_n_shi0 = shr_mem_8_shr_mem_8_or_cse_pff;
  assign din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_8_cns_S0 = ~((shr_mem_8_cns_ppown==2'b10));
  assign shr_mem_8_cns_S0_pff = ~((shr_mem_8_acc_rmff==2'b10));
  assign shr_mem_8_mux_6_nl = MUX_s_1_2_2(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_8_and_3_cse_pff);
  assign shr_mem_8_shr_mem_8_or_cse_pff = (shr_mem_8_mux_6_nl) | (~((shr_mem_8_cns_S0_pff
      & (~ shr_mem_8_xor_rmff)) | shr_mem_8_and_3_cse_pff));
  assign shr_mem_8_cns_csb_n_shi0 = shr_mem_8_shr_mem_8_or_cse_pff;
  assign shr_mem_8_cns_dinb_shi0 = MUX_v_64_2_2(dout_8_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_8_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_8_and_3_cse_pff);
  assign shr_mem_8_cns_addra_shi1 = shr_mem_8_shr_mem_8_mux_2_cse_pff;
  assign shr_mem_8_and_5_cse_pff = shr_mem_8_cns_S1_pff & shr_mem_8_xor_1_rmff;
  assign shr_mem_8_shr_mem_8_mux_2_cse_pff = MUX_v_8_2_2(dout_8_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_8_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_8_and_5_cse_pff);
  assign shr_mem_8_cns_addrb_shi1 = shr_mem_8_shr_mem_8_mux_2_cse_pff;
  assign shr_mem_8_cns_csa_n_shi1 = shr_mem_8_shr_mem_8_or_1_cse_pff;
  assign shr_mem_8_mux_7_nl = MUX_s_1_2_2(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_8_and_5_cse_pff);
  assign shr_mem_8_shr_mem_8_or_1_cse_pff = (shr_mem_8_mux_7_nl) | (~((shr_mem_8_cns_S0_pff
      & shr_mem_8_xor_rmff) | shr_mem_8_and_5_cse_pff));
  assign shr_mem_8_cns_csb_n_shi1 = shr_mem_8_shr_mem_8_or_1_cse_pff;
  assign shr_mem_8_cns_dinb_shi1 = MUX_v_64_2_2(dout_8_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_8_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_8_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_8_cns_ppidx <= 1'b0;
      shr_mem_8_cns_ppown <= 2'b0;
      shr_mem_8_cns_ppidx_1 <= 1'b0;
      shr_mem_8_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_8_cns_ppidx <= shr_mem_8_xor_rmff;
      shr_mem_8_cns_ppown <= shr_mem_8_acc_rmff;
      shr_mem_8_cns_ppidx_1 <= shr_mem_8_xor_1_rmff;
      shr_mem_8_cns_ppown_1 <= shr_mem_8_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeYeetf_7_cns_bctl
// ------------------------------------------------------------------


module double_buffeYeetf_7_cns_bctl (
  clk, rst, dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_7_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_7_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_7_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_7_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_7_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_7_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_7_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_7_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_7_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_7_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_7_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_7_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_7_cns_S0, shr_mem_7_cns_R0, shr_mem_7_cns_S1, shr_mem_7_cns_R1, shr_mem_7_cns_addra_shi0,
      shr_mem_7_cns_addra_shi1, shr_mem_7_cns_addrb_shi0, shr_mem_7_cns_addrb_shi1,
      shr_mem_7_cns_csa_n_shi0, shr_mem_7_cns_csa_n_shi1, shr_mem_7_cns_csb_n_shi0,
      shr_mem_7_cns_csb_n_shi1, shr_mem_7_cns_dinb_shi0, shr_mem_7_cns_dinb_shi1,
      shr_mem_7_cns_douta_sho0, shr_mem_7_cns_douta_sho1, shr_mem_7_cns_S1_pff, din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_7_cns_S0_pff
);
  input clk;
  input rst;
  input dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_7_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_7_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_7_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_7_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_7_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_7_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_7_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_7_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_7_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_7_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_7_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_7_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_7_cns_S0;
  input shr_mem_7_cns_R0;
  output shr_mem_7_cns_S1;
  input shr_mem_7_cns_R1;
  output [7:0] shr_mem_7_cns_addra_shi0;
  output [7:0] shr_mem_7_cns_addra_shi1;
  output [7:0] shr_mem_7_cns_addrb_shi0;
  output [7:0] shr_mem_7_cns_addrb_shi1;
  output shr_mem_7_cns_csa_n_shi0;
  output shr_mem_7_cns_csa_n_shi1;
  output shr_mem_7_cns_csb_n_shi0;
  output shr_mem_7_cns_csb_n_shi1;
  output [63:0] shr_mem_7_cns_dinb_shi0;
  output [63:0] shr_mem_7_cns_dinb_shi1;
  input [63:0] shr_mem_7_cns_douta_sho0;
  input [63:0] shr_mem_7_cns_douta_sho1;
  output shr_mem_7_cns_S1_pff;
  input din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_7_cns_S0_pff;


  // Interconnect Declarations
  reg dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_7_cns_PC0;
  reg shr_mem_7_cns_ppidx;
  reg [1:0] shr_mem_7_cns_ppown;
  wire shr_mem_7_cns_PC1;
  reg shr_mem_7_cns_ppidx_1;
  reg [1:0] shr_mem_7_cns_ppown_1;
  wire [7:0] shr_mem_7_shr_mem_7_mux_3_cse_pff;
  wire shr_mem_7_and_3_cse_pff;
  wire [1:0] shr_mem_7_acc_1_rmff;
  wire [3:0] nl_shr_mem_7_acc_1_rmff;
  wire shr_mem_7_xor_1_rmff;
  wire shr_mem_7_shr_mem_7_or_cse_pff;
  wire [1:0] shr_mem_7_acc_rmff;
  wire [3:0] nl_shr_mem_7_acc_rmff;
  wire shr_mem_7_xor_rmff;
  wire [7:0] shr_mem_7_shr_mem_7_mux_2_cse_pff;
  wire shr_mem_7_and_5_cse_pff;
  wire shr_mem_7_shr_mem_7_or_1_cse_pff;

  wire[0:0] shr_mem_7_mux_6_nl;
  wire[0:0] shr_mem_7_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_7_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_7_cns_R0;
  assign din_7_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_7_cns_R1;
  assign shr_mem_7_xor_rmff = shr_mem_7_cns_ppidx ^ shr_mem_7_cns_PC0;
  assign nl_shr_mem_7_acc_rmff = shr_mem_7_cns_ppown + conv_u2u_1_2(shr_mem_7_cns_PC0)
      + conv_s2u_1_2(shr_mem_7_cns_PC1);
  assign shr_mem_7_acc_rmff = nl_shr_mem_7_acc_rmff[1:0];
  assign shr_mem_7_cns_PC0 = shr_mem_7_cns_S0 & dout_7_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_7_xor_1_rmff = shr_mem_7_cns_ppidx_1 ^ shr_mem_7_cns_PC1;
  assign nl_shr_mem_7_acc_1_rmff = shr_mem_7_cns_ppown_1 + conv_u2u_1_2(shr_mem_7_cns_PC1)
      + conv_s2u_1_2(shr_mem_7_cns_PC0);
  assign shr_mem_7_acc_1_rmff = nl_shr_mem_7_acc_1_rmff[1:0];
  assign shr_mem_7_cns_PC1 = shr_mem_7_cns_S1 & din_7_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_7_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_7_cns_douta_sho0,
      shr_mem_7_cns_douta_sho1, shr_mem_7_cns_ppidx);
  assign din_7_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_7_cns_douta_sho0,
      shr_mem_7_cns_douta_sho1, shr_mem_7_cns_ppidx_1);
  assign shr_mem_7_cns_addra_shi0 = shr_mem_7_shr_mem_7_mux_3_cse_pff;
  assign shr_mem_7_cns_S1 = (shr_mem_7_cns_ppown_1!=2'b00);
  assign shr_mem_7_cns_S1_pff = (shr_mem_7_acc_1_rmff!=2'b00);
  assign shr_mem_7_and_3_cse_pff = shr_mem_7_cns_S1_pff & (~ shr_mem_7_xor_1_rmff);
  assign shr_mem_7_shr_mem_7_mux_3_cse_pff = MUX_v_8_2_2(dout_7_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_7_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_7_and_3_cse_pff);
  assign shr_mem_7_cns_addrb_shi0 = shr_mem_7_shr_mem_7_mux_3_cse_pff;
  assign shr_mem_7_cns_csa_n_shi0 = shr_mem_7_shr_mem_7_or_cse_pff;
  assign din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_7_cns_S0 = ~((shr_mem_7_cns_ppown==2'b10));
  assign shr_mem_7_cns_S0_pff = ~((shr_mem_7_acc_rmff==2'b10));
  assign shr_mem_7_mux_6_nl = MUX_s_1_2_2(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_7_and_3_cse_pff);
  assign shr_mem_7_shr_mem_7_or_cse_pff = (shr_mem_7_mux_6_nl) | (~((shr_mem_7_cns_S0_pff
      & (~ shr_mem_7_xor_rmff)) | shr_mem_7_and_3_cse_pff));
  assign shr_mem_7_cns_csb_n_shi0 = shr_mem_7_shr_mem_7_or_cse_pff;
  assign shr_mem_7_cns_dinb_shi0 = MUX_v_64_2_2(dout_7_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_7_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_7_and_3_cse_pff);
  assign shr_mem_7_cns_addra_shi1 = shr_mem_7_shr_mem_7_mux_2_cse_pff;
  assign shr_mem_7_and_5_cse_pff = shr_mem_7_cns_S1_pff & shr_mem_7_xor_1_rmff;
  assign shr_mem_7_shr_mem_7_mux_2_cse_pff = MUX_v_8_2_2(dout_7_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_7_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_7_and_5_cse_pff);
  assign shr_mem_7_cns_addrb_shi1 = shr_mem_7_shr_mem_7_mux_2_cse_pff;
  assign shr_mem_7_cns_csa_n_shi1 = shr_mem_7_shr_mem_7_or_1_cse_pff;
  assign shr_mem_7_mux_7_nl = MUX_s_1_2_2(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_7_and_5_cse_pff);
  assign shr_mem_7_shr_mem_7_or_1_cse_pff = (shr_mem_7_mux_7_nl) | (~((shr_mem_7_cns_S0_pff
      & shr_mem_7_xor_rmff) | shr_mem_7_and_5_cse_pff));
  assign shr_mem_7_cns_csb_n_shi1 = shr_mem_7_shr_mem_7_or_1_cse_pff;
  assign shr_mem_7_cns_dinb_shi1 = MUX_v_64_2_2(dout_7_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_7_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_7_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_7_cns_ppidx <= 1'b0;
      shr_mem_7_cns_ppown <= 2'b0;
      shr_mem_7_cns_ppidx_1 <= 1'b0;
      shr_mem_7_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_7_cns_ppidx <= shr_mem_7_xor_rmff;
      shr_mem_7_cns_ppown <= shr_mem_7_acc_rmff;
      shr_mem_7_cns_ppidx_1 <= shr_mem_7_xor_1_rmff;
      shr_mem_7_cns_ppown_1 <= shr_mem_7_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeYeetf_6_cns_bctl
// ------------------------------------------------------------------


module double_buffeYeetf_6_cns_bctl (
  clk, rst, dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_6_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_6_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_6_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_6_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_6_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_6_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_6_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_6_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_6_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_6_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_6_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_6_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_6_cns_S0, shr_mem_6_cns_R0, shr_mem_6_cns_S1, shr_mem_6_cns_R1, shr_mem_6_cns_addra_shi0,
      shr_mem_6_cns_addra_shi1, shr_mem_6_cns_addrb_shi0, shr_mem_6_cns_addrb_shi1,
      shr_mem_6_cns_csa_n_shi0, shr_mem_6_cns_csa_n_shi1, shr_mem_6_cns_csb_n_shi0,
      shr_mem_6_cns_csb_n_shi1, shr_mem_6_cns_dinb_shi0, shr_mem_6_cns_dinb_shi1,
      shr_mem_6_cns_douta_sho0, shr_mem_6_cns_douta_sho1, shr_mem_6_cns_S1_pff, din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_6_cns_S0_pff
);
  input clk;
  input rst;
  input dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_6_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_6_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_6_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_6_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_6_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_6_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_6_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_6_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_6_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_6_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_6_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_6_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_6_cns_S0;
  input shr_mem_6_cns_R0;
  output shr_mem_6_cns_S1;
  input shr_mem_6_cns_R1;
  output [7:0] shr_mem_6_cns_addra_shi0;
  output [7:0] shr_mem_6_cns_addra_shi1;
  output [7:0] shr_mem_6_cns_addrb_shi0;
  output [7:0] shr_mem_6_cns_addrb_shi1;
  output shr_mem_6_cns_csa_n_shi0;
  output shr_mem_6_cns_csa_n_shi1;
  output shr_mem_6_cns_csb_n_shi0;
  output shr_mem_6_cns_csb_n_shi1;
  output [63:0] shr_mem_6_cns_dinb_shi0;
  output [63:0] shr_mem_6_cns_dinb_shi1;
  input [63:0] shr_mem_6_cns_douta_sho0;
  input [63:0] shr_mem_6_cns_douta_sho1;
  output shr_mem_6_cns_S1_pff;
  input din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_6_cns_S0_pff;


  // Interconnect Declarations
  reg dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_6_cns_PC0;
  reg shr_mem_6_cns_ppidx;
  reg [1:0] shr_mem_6_cns_ppown;
  wire shr_mem_6_cns_PC1;
  reg shr_mem_6_cns_ppidx_1;
  reg [1:0] shr_mem_6_cns_ppown_1;
  wire [7:0] shr_mem_6_shr_mem_6_mux_3_cse_pff;
  wire shr_mem_6_and_3_cse_pff;
  wire [1:0] shr_mem_6_acc_1_rmff;
  wire [3:0] nl_shr_mem_6_acc_1_rmff;
  wire shr_mem_6_xor_1_rmff;
  wire shr_mem_6_shr_mem_6_or_cse_pff;
  wire [1:0] shr_mem_6_acc_rmff;
  wire [3:0] nl_shr_mem_6_acc_rmff;
  wire shr_mem_6_xor_rmff;
  wire [7:0] shr_mem_6_shr_mem_6_mux_2_cse_pff;
  wire shr_mem_6_and_5_cse_pff;
  wire shr_mem_6_shr_mem_6_or_1_cse_pff;

  wire[0:0] shr_mem_6_mux_6_nl;
  wire[0:0] shr_mem_6_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_6_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_6_cns_R0;
  assign din_6_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_6_cns_R1;
  assign shr_mem_6_xor_rmff = shr_mem_6_cns_ppidx ^ shr_mem_6_cns_PC0;
  assign nl_shr_mem_6_acc_rmff = shr_mem_6_cns_ppown + conv_u2u_1_2(shr_mem_6_cns_PC0)
      + conv_s2u_1_2(shr_mem_6_cns_PC1);
  assign shr_mem_6_acc_rmff = nl_shr_mem_6_acc_rmff[1:0];
  assign shr_mem_6_cns_PC0 = shr_mem_6_cns_S0 & dout_6_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_6_xor_1_rmff = shr_mem_6_cns_ppidx_1 ^ shr_mem_6_cns_PC1;
  assign nl_shr_mem_6_acc_1_rmff = shr_mem_6_cns_ppown_1 + conv_u2u_1_2(shr_mem_6_cns_PC1)
      + conv_s2u_1_2(shr_mem_6_cns_PC0);
  assign shr_mem_6_acc_1_rmff = nl_shr_mem_6_acc_1_rmff[1:0];
  assign shr_mem_6_cns_PC1 = shr_mem_6_cns_S1 & din_6_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_6_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_6_cns_douta_sho0,
      shr_mem_6_cns_douta_sho1, shr_mem_6_cns_ppidx);
  assign din_6_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_6_cns_douta_sho0,
      shr_mem_6_cns_douta_sho1, shr_mem_6_cns_ppidx_1);
  assign shr_mem_6_cns_addra_shi0 = shr_mem_6_shr_mem_6_mux_3_cse_pff;
  assign shr_mem_6_cns_S1 = (shr_mem_6_cns_ppown_1!=2'b00);
  assign shr_mem_6_cns_S1_pff = (shr_mem_6_acc_1_rmff!=2'b00);
  assign shr_mem_6_and_3_cse_pff = shr_mem_6_cns_S1_pff & (~ shr_mem_6_xor_1_rmff);
  assign shr_mem_6_shr_mem_6_mux_3_cse_pff = MUX_v_8_2_2(dout_6_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_6_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_6_and_3_cse_pff);
  assign shr_mem_6_cns_addrb_shi0 = shr_mem_6_shr_mem_6_mux_3_cse_pff;
  assign shr_mem_6_cns_csa_n_shi0 = shr_mem_6_shr_mem_6_or_cse_pff;
  assign din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_6_cns_S0 = ~((shr_mem_6_cns_ppown==2'b10));
  assign shr_mem_6_cns_S0_pff = ~((shr_mem_6_acc_rmff==2'b10));
  assign shr_mem_6_mux_6_nl = MUX_s_1_2_2(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_6_and_3_cse_pff);
  assign shr_mem_6_shr_mem_6_or_cse_pff = (shr_mem_6_mux_6_nl) | (~((shr_mem_6_cns_S0_pff
      & (~ shr_mem_6_xor_rmff)) | shr_mem_6_and_3_cse_pff));
  assign shr_mem_6_cns_csb_n_shi0 = shr_mem_6_shr_mem_6_or_cse_pff;
  assign shr_mem_6_cns_dinb_shi0 = MUX_v_64_2_2(dout_6_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_6_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_6_and_3_cse_pff);
  assign shr_mem_6_cns_addra_shi1 = shr_mem_6_shr_mem_6_mux_2_cse_pff;
  assign shr_mem_6_and_5_cse_pff = shr_mem_6_cns_S1_pff & shr_mem_6_xor_1_rmff;
  assign shr_mem_6_shr_mem_6_mux_2_cse_pff = MUX_v_8_2_2(dout_6_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_6_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_6_and_5_cse_pff);
  assign shr_mem_6_cns_addrb_shi1 = shr_mem_6_shr_mem_6_mux_2_cse_pff;
  assign shr_mem_6_cns_csa_n_shi1 = shr_mem_6_shr_mem_6_or_1_cse_pff;
  assign shr_mem_6_mux_7_nl = MUX_s_1_2_2(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_6_and_5_cse_pff);
  assign shr_mem_6_shr_mem_6_or_1_cse_pff = (shr_mem_6_mux_7_nl) | (~((shr_mem_6_cns_S0_pff
      & shr_mem_6_xor_rmff) | shr_mem_6_and_5_cse_pff));
  assign shr_mem_6_cns_csb_n_shi1 = shr_mem_6_shr_mem_6_or_1_cse_pff;
  assign shr_mem_6_cns_dinb_shi1 = MUX_v_64_2_2(dout_6_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_6_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_6_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_6_cns_ppidx <= 1'b0;
      shr_mem_6_cns_ppown <= 2'b0;
      shr_mem_6_cns_ppidx_1 <= 1'b0;
      shr_mem_6_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_6_cns_ppidx <= shr_mem_6_xor_rmff;
      shr_mem_6_cns_ppown <= shr_mem_6_acc_rmff;
      shr_mem_6_cns_ppidx_1 <= shr_mem_6_xor_1_rmff;
      shr_mem_6_cns_ppown_1 <= shr_mem_6_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeYeetf_5_cns_bctl
// ------------------------------------------------------------------


module double_buffeYeetf_5_cns_bctl (
  clk, rst, dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_5_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_5_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_5_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_5_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_5_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_5_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_5_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_5_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_5_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_5_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_5_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_5_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_5_cns_S0, shr_mem_5_cns_R0, shr_mem_5_cns_S1, shr_mem_5_cns_R1, shr_mem_5_cns_addra_shi0,
      shr_mem_5_cns_addra_shi1, shr_mem_5_cns_addrb_shi0, shr_mem_5_cns_addrb_shi1,
      shr_mem_5_cns_csa_n_shi0, shr_mem_5_cns_csa_n_shi1, shr_mem_5_cns_csb_n_shi0,
      shr_mem_5_cns_csb_n_shi1, shr_mem_5_cns_dinb_shi0, shr_mem_5_cns_dinb_shi1,
      shr_mem_5_cns_douta_sho0, shr_mem_5_cns_douta_sho1, shr_mem_5_cns_S1_pff, din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_5_cns_S0_pff
);
  input clk;
  input rst;
  input dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_5_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_5_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_5_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_5_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_5_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_5_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_5_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_5_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_5_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_5_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_5_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_5_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_5_cns_S0;
  input shr_mem_5_cns_R0;
  output shr_mem_5_cns_S1;
  input shr_mem_5_cns_R1;
  output [7:0] shr_mem_5_cns_addra_shi0;
  output [7:0] shr_mem_5_cns_addra_shi1;
  output [7:0] shr_mem_5_cns_addrb_shi0;
  output [7:0] shr_mem_5_cns_addrb_shi1;
  output shr_mem_5_cns_csa_n_shi0;
  output shr_mem_5_cns_csa_n_shi1;
  output shr_mem_5_cns_csb_n_shi0;
  output shr_mem_5_cns_csb_n_shi1;
  output [63:0] shr_mem_5_cns_dinb_shi0;
  output [63:0] shr_mem_5_cns_dinb_shi1;
  input [63:0] shr_mem_5_cns_douta_sho0;
  input [63:0] shr_mem_5_cns_douta_sho1;
  output shr_mem_5_cns_S1_pff;
  input din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_5_cns_S0_pff;


  // Interconnect Declarations
  reg dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_5_cns_PC0;
  reg shr_mem_5_cns_ppidx;
  reg [1:0] shr_mem_5_cns_ppown;
  wire shr_mem_5_cns_PC1;
  reg shr_mem_5_cns_ppidx_1;
  reg [1:0] shr_mem_5_cns_ppown_1;
  wire [7:0] shr_mem_5_shr_mem_5_mux_3_cse_pff;
  wire shr_mem_5_and_3_cse_pff;
  wire [1:0] shr_mem_5_acc_1_rmff;
  wire [3:0] nl_shr_mem_5_acc_1_rmff;
  wire shr_mem_5_xor_1_rmff;
  wire shr_mem_5_shr_mem_5_or_cse_pff;
  wire [1:0] shr_mem_5_acc_rmff;
  wire [3:0] nl_shr_mem_5_acc_rmff;
  wire shr_mem_5_xor_rmff;
  wire [7:0] shr_mem_5_shr_mem_5_mux_2_cse_pff;
  wire shr_mem_5_and_5_cse_pff;
  wire shr_mem_5_shr_mem_5_or_1_cse_pff;

  wire[0:0] shr_mem_5_mux_6_nl;
  wire[0:0] shr_mem_5_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_5_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_5_cns_R0;
  assign din_5_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_5_cns_R1;
  assign shr_mem_5_xor_rmff = shr_mem_5_cns_ppidx ^ shr_mem_5_cns_PC0;
  assign nl_shr_mem_5_acc_rmff = shr_mem_5_cns_ppown + conv_u2u_1_2(shr_mem_5_cns_PC0)
      + conv_s2u_1_2(shr_mem_5_cns_PC1);
  assign shr_mem_5_acc_rmff = nl_shr_mem_5_acc_rmff[1:0];
  assign shr_mem_5_cns_PC0 = shr_mem_5_cns_S0 & dout_5_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_5_xor_1_rmff = shr_mem_5_cns_ppidx_1 ^ shr_mem_5_cns_PC1;
  assign nl_shr_mem_5_acc_1_rmff = shr_mem_5_cns_ppown_1 + conv_u2u_1_2(shr_mem_5_cns_PC1)
      + conv_s2u_1_2(shr_mem_5_cns_PC0);
  assign shr_mem_5_acc_1_rmff = nl_shr_mem_5_acc_1_rmff[1:0];
  assign shr_mem_5_cns_PC1 = shr_mem_5_cns_S1 & din_5_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_5_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_5_cns_douta_sho0,
      shr_mem_5_cns_douta_sho1, shr_mem_5_cns_ppidx);
  assign din_5_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_5_cns_douta_sho0,
      shr_mem_5_cns_douta_sho1, shr_mem_5_cns_ppidx_1);
  assign shr_mem_5_cns_addra_shi0 = shr_mem_5_shr_mem_5_mux_3_cse_pff;
  assign shr_mem_5_cns_S1 = (shr_mem_5_cns_ppown_1!=2'b00);
  assign shr_mem_5_cns_S1_pff = (shr_mem_5_acc_1_rmff!=2'b00);
  assign shr_mem_5_and_3_cse_pff = shr_mem_5_cns_S1_pff & (~ shr_mem_5_xor_1_rmff);
  assign shr_mem_5_shr_mem_5_mux_3_cse_pff = MUX_v_8_2_2(dout_5_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_5_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_5_and_3_cse_pff);
  assign shr_mem_5_cns_addrb_shi0 = shr_mem_5_shr_mem_5_mux_3_cse_pff;
  assign shr_mem_5_cns_csa_n_shi0 = shr_mem_5_shr_mem_5_or_cse_pff;
  assign din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_5_cns_S0 = ~((shr_mem_5_cns_ppown==2'b10));
  assign shr_mem_5_cns_S0_pff = ~((shr_mem_5_acc_rmff==2'b10));
  assign shr_mem_5_mux_6_nl = MUX_s_1_2_2(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_5_and_3_cse_pff);
  assign shr_mem_5_shr_mem_5_or_cse_pff = (shr_mem_5_mux_6_nl) | (~((shr_mem_5_cns_S0_pff
      & (~ shr_mem_5_xor_rmff)) | shr_mem_5_and_3_cse_pff));
  assign shr_mem_5_cns_csb_n_shi0 = shr_mem_5_shr_mem_5_or_cse_pff;
  assign shr_mem_5_cns_dinb_shi0 = MUX_v_64_2_2(dout_5_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_5_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_5_and_3_cse_pff);
  assign shr_mem_5_cns_addra_shi1 = shr_mem_5_shr_mem_5_mux_2_cse_pff;
  assign shr_mem_5_and_5_cse_pff = shr_mem_5_cns_S1_pff & shr_mem_5_xor_1_rmff;
  assign shr_mem_5_shr_mem_5_mux_2_cse_pff = MUX_v_8_2_2(dout_5_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_5_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_5_and_5_cse_pff);
  assign shr_mem_5_cns_addrb_shi1 = shr_mem_5_shr_mem_5_mux_2_cse_pff;
  assign shr_mem_5_cns_csa_n_shi1 = shr_mem_5_shr_mem_5_or_1_cse_pff;
  assign shr_mem_5_mux_7_nl = MUX_s_1_2_2(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_5_and_5_cse_pff);
  assign shr_mem_5_shr_mem_5_or_1_cse_pff = (shr_mem_5_mux_7_nl) | (~((shr_mem_5_cns_S0_pff
      & shr_mem_5_xor_rmff) | shr_mem_5_and_5_cse_pff));
  assign shr_mem_5_cns_csb_n_shi1 = shr_mem_5_shr_mem_5_or_1_cse_pff;
  assign shr_mem_5_cns_dinb_shi1 = MUX_v_64_2_2(dout_5_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_5_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_5_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_5_cns_ppidx <= 1'b0;
      shr_mem_5_cns_ppown <= 2'b0;
      shr_mem_5_cns_ppidx_1 <= 1'b0;
      shr_mem_5_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_5_cns_ppidx <= shr_mem_5_xor_rmff;
      shr_mem_5_cns_ppown <= shr_mem_5_acc_rmff;
      shr_mem_5_cns_ppidx_1 <= shr_mem_5_xor_1_rmff;
      shr_mem_5_cns_ppown_1 <= shr_mem_5_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeYeetf_4_cns_bctl
// ------------------------------------------------------------------


module double_buffeYeetf_4_cns_bctl (
  clk, rst, dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_4_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_4_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_4_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_4_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_4_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_4_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_4_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_4_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_4_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_4_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_4_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_4_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_4_cns_S0, shr_mem_4_cns_R0, shr_mem_4_cns_S1, shr_mem_4_cns_R1, shr_mem_4_cns_addra_shi0,
      shr_mem_4_cns_addra_shi1, shr_mem_4_cns_addrb_shi0, shr_mem_4_cns_addrb_shi1,
      shr_mem_4_cns_csa_n_shi0, shr_mem_4_cns_csa_n_shi1, shr_mem_4_cns_csb_n_shi0,
      shr_mem_4_cns_csb_n_shi1, shr_mem_4_cns_dinb_shi0, shr_mem_4_cns_dinb_shi1,
      shr_mem_4_cns_douta_sho0, shr_mem_4_cns_douta_sho1, shr_mem_4_cns_S1_pff, din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_4_cns_S0_pff
);
  input clk;
  input rst;
  input dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_4_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_4_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_4_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_4_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_4_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_4_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_4_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_4_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_4_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_4_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_4_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_4_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_4_cns_S0;
  input shr_mem_4_cns_R0;
  output shr_mem_4_cns_S1;
  input shr_mem_4_cns_R1;
  output [7:0] shr_mem_4_cns_addra_shi0;
  output [7:0] shr_mem_4_cns_addra_shi1;
  output [7:0] shr_mem_4_cns_addrb_shi0;
  output [7:0] shr_mem_4_cns_addrb_shi1;
  output shr_mem_4_cns_csa_n_shi0;
  output shr_mem_4_cns_csa_n_shi1;
  output shr_mem_4_cns_csb_n_shi0;
  output shr_mem_4_cns_csb_n_shi1;
  output [63:0] shr_mem_4_cns_dinb_shi0;
  output [63:0] shr_mem_4_cns_dinb_shi1;
  input [63:0] shr_mem_4_cns_douta_sho0;
  input [63:0] shr_mem_4_cns_douta_sho1;
  output shr_mem_4_cns_S1_pff;
  input din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_4_cns_S0_pff;


  // Interconnect Declarations
  reg dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_4_cns_PC0;
  reg shr_mem_4_cns_ppidx;
  reg [1:0] shr_mem_4_cns_ppown;
  wire shr_mem_4_cns_PC1;
  reg shr_mem_4_cns_ppidx_1;
  reg [1:0] shr_mem_4_cns_ppown_1;
  wire [7:0] shr_mem_4_shr_mem_4_mux_3_cse_pff;
  wire shr_mem_4_and_3_cse_pff;
  wire [1:0] shr_mem_4_acc_1_rmff;
  wire [3:0] nl_shr_mem_4_acc_1_rmff;
  wire shr_mem_4_xor_1_rmff;
  wire shr_mem_4_shr_mem_4_or_cse_pff;
  wire [1:0] shr_mem_4_acc_rmff;
  wire [3:0] nl_shr_mem_4_acc_rmff;
  wire shr_mem_4_xor_rmff;
  wire [7:0] shr_mem_4_shr_mem_4_mux_2_cse_pff;
  wire shr_mem_4_and_5_cse_pff;
  wire shr_mem_4_shr_mem_4_or_1_cse_pff;

  wire[0:0] shr_mem_4_mux_6_nl;
  wire[0:0] shr_mem_4_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_4_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_4_cns_R0;
  assign din_4_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_4_cns_R1;
  assign shr_mem_4_xor_rmff = shr_mem_4_cns_ppidx ^ shr_mem_4_cns_PC0;
  assign nl_shr_mem_4_acc_rmff = shr_mem_4_cns_ppown + conv_u2u_1_2(shr_mem_4_cns_PC0)
      + conv_s2u_1_2(shr_mem_4_cns_PC1);
  assign shr_mem_4_acc_rmff = nl_shr_mem_4_acc_rmff[1:0];
  assign shr_mem_4_cns_PC0 = shr_mem_4_cns_S0 & dout_4_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_4_xor_1_rmff = shr_mem_4_cns_ppidx_1 ^ shr_mem_4_cns_PC1;
  assign nl_shr_mem_4_acc_1_rmff = shr_mem_4_cns_ppown_1 + conv_u2u_1_2(shr_mem_4_cns_PC1)
      + conv_s2u_1_2(shr_mem_4_cns_PC0);
  assign shr_mem_4_acc_1_rmff = nl_shr_mem_4_acc_1_rmff[1:0];
  assign shr_mem_4_cns_PC1 = shr_mem_4_cns_S1 & din_4_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_4_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_4_cns_douta_sho0,
      shr_mem_4_cns_douta_sho1, shr_mem_4_cns_ppidx);
  assign din_4_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_4_cns_douta_sho0,
      shr_mem_4_cns_douta_sho1, shr_mem_4_cns_ppidx_1);
  assign shr_mem_4_cns_addra_shi0 = shr_mem_4_shr_mem_4_mux_3_cse_pff;
  assign shr_mem_4_cns_S1 = (shr_mem_4_cns_ppown_1!=2'b00);
  assign shr_mem_4_cns_S1_pff = (shr_mem_4_acc_1_rmff!=2'b00);
  assign shr_mem_4_and_3_cse_pff = shr_mem_4_cns_S1_pff & (~ shr_mem_4_xor_1_rmff);
  assign shr_mem_4_shr_mem_4_mux_3_cse_pff = MUX_v_8_2_2(dout_4_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_4_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_4_and_3_cse_pff);
  assign shr_mem_4_cns_addrb_shi0 = shr_mem_4_shr_mem_4_mux_3_cse_pff;
  assign shr_mem_4_cns_csa_n_shi0 = shr_mem_4_shr_mem_4_or_cse_pff;
  assign din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_4_cns_S0 = ~((shr_mem_4_cns_ppown==2'b10));
  assign shr_mem_4_cns_S0_pff = ~((shr_mem_4_acc_rmff==2'b10));
  assign shr_mem_4_mux_6_nl = MUX_s_1_2_2(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_4_and_3_cse_pff);
  assign shr_mem_4_shr_mem_4_or_cse_pff = (shr_mem_4_mux_6_nl) | (~((shr_mem_4_cns_S0_pff
      & (~ shr_mem_4_xor_rmff)) | shr_mem_4_and_3_cse_pff));
  assign shr_mem_4_cns_csb_n_shi0 = shr_mem_4_shr_mem_4_or_cse_pff;
  assign shr_mem_4_cns_dinb_shi0 = MUX_v_64_2_2(dout_4_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_4_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_4_and_3_cse_pff);
  assign shr_mem_4_cns_addra_shi1 = shr_mem_4_shr_mem_4_mux_2_cse_pff;
  assign shr_mem_4_and_5_cse_pff = shr_mem_4_cns_S1_pff & shr_mem_4_xor_1_rmff;
  assign shr_mem_4_shr_mem_4_mux_2_cse_pff = MUX_v_8_2_2(dout_4_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_4_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_4_and_5_cse_pff);
  assign shr_mem_4_cns_addrb_shi1 = shr_mem_4_shr_mem_4_mux_2_cse_pff;
  assign shr_mem_4_cns_csa_n_shi1 = shr_mem_4_shr_mem_4_or_1_cse_pff;
  assign shr_mem_4_mux_7_nl = MUX_s_1_2_2(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_4_and_5_cse_pff);
  assign shr_mem_4_shr_mem_4_or_1_cse_pff = (shr_mem_4_mux_7_nl) | (~((shr_mem_4_cns_S0_pff
      & shr_mem_4_xor_rmff) | shr_mem_4_and_5_cse_pff));
  assign shr_mem_4_cns_csb_n_shi1 = shr_mem_4_shr_mem_4_or_1_cse_pff;
  assign shr_mem_4_cns_dinb_shi1 = MUX_v_64_2_2(dout_4_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_4_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_4_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_4_cns_ppidx <= 1'b0;
      shr_mem_4_cns_ppown <= 2'b0;
      shr_mem_4_cns_ppidx_1 <= 1'b0;
      shr_mem_4_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_4_cns_ppidx <= shr_mem_4_xor_rmff;
      shr_mem_4_cns_ppown <= shr_mem_4_acc_rmff;
      shr_mem_4_cns_ppidx_1 <= shr_mem_4_xor_1_rmff;
      shr_mem_4_cns_ppown_1 <= shr_mem_4_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeYeetf_3_cns_bctl
// ------------------------------------------------------------------


module double_buffeYeetf_3_cns_bctl (
  clk, rst, dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_3_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_3_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_3_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_3_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_3_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_3_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_3_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_3_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_3_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_3_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_3_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_3_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_3_cns_S0, shr_mem_3_cns_R0, shr_mem_3_cns_S1, shr_mem_3_cns_R1, shr_mem_3_cns_addra_shi0,
      shr_mem_3_cns_addra_shi1, shr_mem_3_cns_addrb_shi0, shr_mem_3_cns_addrb_shi1,
      shr_mem_3_cns_csa_n_shi0, shr_mem_3_cns_csa_n_shi1, shr_mem_3_cns_csb_n_shi0,
      shr_mem_3_cns_csb_n_shi1, shr_mem_3_cns_dinb_shi0, shr_mem_3_cns_dinb_shi1,
      shr_mem_3_cns_douta_sho0, shr_mem_3_cns_douta_sho1, shr_mem_3_cns_S1_pff, din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_3_cns_S0_pff
);
  input clk;
  input rst;
  input dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_3_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_3_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_3_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_3_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_3_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_3_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_3_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_3_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_3_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_3_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_3_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_3_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_3_cns_S0;
  input shr_mem_3_cns_R0;
  output shr_mem_3_cns_S1;
  input shr_mem_3_cns_R1;
  output [7:0] shr_mem_3_cns_addra_shi0;
  output [7:0] shr_mem_3_cns_addra_shi1;
  output [7:0] shr_mem_3_cns_addrb_shi0;
  output [7:0] shr_mem_3_cns_addrb_shi1;
  output shr_mem_3_cns_csa_n_shi0;
  output shr_mem_3_cns_csa_n_shi1;
  output shr_mem_3_cns_csb_n_shi0;
  output shr_mem_3_cns_csb_n_shi1;
  output [63:0] shr_mem_3_cns_dinb_shi0;
  output [63:0] shr_mem_3_cns_dinb_shi1;
  input [63:0] shr_mem_3_cns_douta_sho0;
  input [63:0] shr_mem_3_cns_douta_sho1;
  output shr_mem_3_cns_S1_pff;
  input din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_3_cns_S0_pff;


  // Interconnect Declarations
  reg dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_3_cns_PC0;
  reg shr_mem_3_cns_ppidx;
  reg [1:0] shr_mem_3_cns_ppown;
  wire shr_mem_3_cns_PC1;
  reg shr_mem_3_cns_ppidx_1;
  reg [1:0] shr_mem_3_cns_ppown_1;
  wire [7:0] shr_mem_3_shr_mem_3_mux_3_cse_pff;
  wire shr_mem_3_and_3_cse_pff;
  wire [1:0] shr_mem_3_acc_1_rmff;
  wire [3:0] nl_shr_mem_3_acc_1_rmff;
  wire shr_mem_3_xor_1_rmff;
  wire shr_mem_3_shr_mem_3_or_cse_pff;
  wire [1:0] shr_mem_3_acc_rmff;
  wire [3:0] nl_shr_mem_3_acc_rmff;
  wire shr_mem_3_xor_rmff;
  wire [7:0] shr_mem_3_shr_mem_3_mux_2_cse_pff;
  wire shr_mem_3_and_5_cse_pff;
  wire shr_mem_3_shr_mem_3_or_1_cse_pff;

  wire[0:0] shr_mem_3_mux_6_nl;
  wire[0:0] shr_mem_3_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_3_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_3_cns_R0;
  assign din_3_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_3_cns_R1;
  assign shr_mem_3_xor_rmff = shr_mem_3_cns_ppidx ^ shr_mem_3_cns_PC0;
  assign nl_shr_mem_3_acc_rmff = shr_mem_3_cns_ppown + conv_u2u_1_2(shr_mem_3_cns_PC0)
      + conv_s2u_1_2(shr_mem_3_cns_PC1);
  assign shr_mem_3_acc_rmff = nl_shr_mem_3_acc_rmff[1:0];
  assign shr_mem_3_cns_PC0 = shr_mem_3_cns_S0 & dout_3_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_3_xor_1_rmff = shr_mem_3_cns_ppidx_1 ^ shr_mem_3_cns_PC1;
  assign nl_shr_mem_3_acc_1_rmff = shr_mem_3_cns_ppown_1 + conv_u2u_1_2(shr_mem_3_cns_PC1)
      + conv_s2u_1_2(shr_mem_3_cns_PC0);
  assign shr_mem_3_acc_1_rmff = nl_shr_mem_3_acc_1_rmff[1:0];
  assign shr_mem_3_cns_PC1 = shr_mem_3_cns_S1 & din_3_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_3_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_3_cns_douta_sho0,
      shr_mem_3_cns_douta_sho1, shr_mem_3_cns_ppidx);
  assign din_3_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_3_cns_douta_sho0,
      shr_mem_3_cns_douta_sho1, shr_mem_3_cns_ppidx_1);
  assign shr_mem_3_cns_addra_shi0 = shr_mem_3_shr_mem_3_mux_3_cse_pff;
  assign shr_mem_3_cns_S1 = (shr_mem_3_cns_ppown_1!=2'b00);
  assign shr_mem_3_cns_S1_pff = (shr_mem_3_acc_1_rmff!=2'b00);
  assign shr_mem_3_and_3_cse_pff = shr_mem_3_cns_S1_pff & (~ shr_mem_3_xor_1_rmff);
  assign shr_mem_3_shr_mem_3_mux_3_cse_pff = MUX_v_8_2_2(dout_3_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_3_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_3_and_3_cse_pff);
  assign shr_mem_3_cns_addrb_shi0 = shr_mem_3_shr_mem_3_mux_3_cse_pff;
  assign shr_mem_3_cns_csa_n_shi0 = shr_mem_3_shr_mem_3_or_cse_pff;
  assign din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_3_cns_S0 = ~((shr_mem_3_cns_ppown==2'b10));
  assign shr_mem_3_cns_S0_pff = ~((shr_mem_3_acc_rmff==2'b10));
  assign shr_mem_3_mux_6_nl = MUX_s_1_2_2(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_3_and_3_cse_pff);
  assign shr_mem_3_shr_mem_3_or_cse_pff = (shr_mem_3_mux_6_nl) | (~((shr_mem_3_cns_S0_pff
      & (~ shr_mem_3_xor_rmff)) | shr_mem_3_and_3_cse_pff));
  assign shr_mem_3_cns_csb_n_shi0 = shr_mem_3_shr_mem_3_or_cse_pff;
  assign shr_mem_3_cns_dinb_shi0 = MUX_v_64_2_2(dout_3_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_3_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_3_and_3_cse_pff);
  assign shr_mem_3_cns_addra_shi1 = shr_mem_3_shr_mem_3_mux_2_cse_pff;
  assign shr_mem_3_and_5_cse_pff = shr_mem_3_cns_S1_pff & shr_mem_3_xor_1_rmff;
  assign shr_mem_3_shr_mem_3_mux_2_cse_pff = MUX_v_8_2_2(dout_3_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_3_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_3_and_5_cse_pff);
  assign shr_mem_3_cns_addrb_shi1 = shr_mem_3_shr_mem_3_mux_2_cse_pff;
  assign shr_mem_3_cns_csa_n_shi1 = shr_mem_3_shr_mem_3_or_1_cse_pff;
  assign shr_mem_3_mux_7_nl = MUX_s_1_2_2(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_3_and_5_cse_pff);
  assign shr_mem_3_shr_mem_3_or_1_cse_pff = (shr_mem_3_mux_7_nl) | (~((shr_mem_3_cns_S0_pff
      & shr_mem_3_xor_rmff) | shr_mem_3_and_5_cse_pff));
  assign shr_mem_3_cns_csb_n_shi1 = shr_mem_3_shr_mem_3_or_1_cse_pff;
  assign shr_mem_3_cns_dinb_shi1 = MUX_v_64_2_2(dout_3_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_3_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_3_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_3_cns_ppidx <= 1'b0;
      shr_mem_3_cns_ppown <= 2'b0;
      shr_mem_3_cns_ppidx_1 <= 1'b0;
      shr_mem_3_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_3_cns_ppidx <= shr_mem_3_xor_rmff;
      shr_mem_3_cns_ppown <= shr_mem_3_acc_rmff;
      shr_mem_3_cns_ppidx_1 <= shr_mem_3_xor_1_rmff;
      shr_mem_3_cns_ppown_1 <= shr_mem_3_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeYeetf_2_cns_bctl
// ------------------------------------------------------------------


module double_buffeYeetf_2_cns_bctl (
  clk, rst, dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_2_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_2_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_2_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_2_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_2_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_2_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_2_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_2_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_2_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_2_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_2_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_2_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_2_cns_S0, shr_mem_2_cns_R0, shr_mem_2_cns_S1, shr_mem_2_cns_R1, shr_mem_2_cns_addra_shi0,
      shr_mem_2_cns_addra_shi1, shr_mem_2_cns_addrb_shi0, shr_mem_2_cns_addrb_shi1,
      shr_mem_2_cns_csa_n_shi0, shr_mem_2_cns_csa_n_shi1, shr_mem_2_cns_csb_n_shi0,
      shr_mem_2_cns_csb_n_shi1, shr_mem_2_cns_dinb_shi0, shr_mem_2_cns_dinb_shi1,
      shr_mem_2_cns_douta_sho0, shr_mem_2_cns_douta_sho1, shr_mem_2_cns_S1_pff, din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_2_cns_S0_pff
);
  input clk;
  input rst;
  input dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_2_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_2_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_2_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_2_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_2_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_2_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_2_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_2_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_2_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_2_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_2_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_2_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_2_cns_S0;
  input shr_mem_2_cns_R0;
  output shr_mem_2_cns_S1;
  input shr_mem_2_cns_R1;
  output [7:0] shr_mem_2_cns_addra_shi0;
  output [7:0] shr_mem_2_cns_addra_shi1;
  output [7:0] shr_mem_2_cns_addrb_shi0;
  output [7:0] shr_mem_2_cns_addrb_shi1;
  output shr_mem_2_cns_csa_n_shi0;
  output shr_mem_2_cns_csa_n_shi1;
  output shr_mem_2_cns_csb_n_shi0;
  output shr_mem_2_cns_csb_n_shi1;
  output [63:0] shr_mem_2_cns_dinb_shi0;
  output [63:0] shr_mem_2_cns_dinb_shi1;
  input [63:0] shr_mem_2_cns_douta_sho0;
  input [63:0] shr_mem_2_cns_douta_sho1;
  output shr_mem_2_cns_S1_pff;
  input din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_2_cns_S0_pff;


  // Interconnect Declarations
  reg dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_2_cns_PC0;
  reg shr_mem_2_cns_ppidx;
  reg [1:0] shr_mem_2_cns_ppown;
  wire shr_mem_2_cns_PC1;
  reg shr_mem_2_cns_ppidx_1;
  reg [1:0] shr_mem_2_cns_ppown_1;
  wire [7:0] shr_mem_2_shr_mem_2_mux_3_cse_pff;
  wire shr_mem_2_and_3_cse_pff;
  wire [1:0] shr_mem_2_acc_1_rmff;
  wire [3:0] nl_shr_mem_2_acc_1_rmff;
  wire shr_mem_2_xor_1_rmff;
  wire shr_mem_2_shr_mem_2_or_cse_pff;
  wire [1:0] shr_mem_2_acc_rmff;
  wire [3:0] nl_shr_mem_2_acc_rmff;
  wire shr_mem_2_xor_rmff;
  wire [7:0] shr_mem_2_shr_mem_2_mux_2_cse_pff;
  wire shr_mem_2_and_5_cse_pff;
  wire shr_mem_2_shr_mem_2_or_1_cse_pff;

  wire[0:0] shr_mem_2_mux_6_nl;
  wire[0:0] shr_mem_2_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_2_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_2_cns_R0;
  assign din_2_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_2_cns_R1;
  assign shr_mem_2_xor_rmff = shr_mem_2_cns_ppidx ^ shr_mem_2_cns_PC0;
  assign nl_shr_mem_2_acc_rmff = shr_mem_2_cns_ppown + conv_u2u_1_2(shr_mem_2_cns_PC0)
      + conv_s2u_1_2(shr_mem_2_cns_PC1);
  assign shr_mem_2_acc_rmff = nl_shr_mem_2_acc_rmff[1:0];
  assign shr_mem_2_cns_PC0 = shr_mem_2_cns_S0 & dout_2_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_2_xor_1_rmff = shr_mem_2_cns_ppidx_1 ^ shr_mem_2_cns_PC1;
  assign nl_shr_mem_2_acc_1_rmff = shr_mem_2_cns_ppown_1 + conv_u2u_1_2(shr_mem_2_cns_PC1)
      + conv_s2u_1_2(shr_mem_2_cns_PC0);
  assign shr_mem_2_acc_1_rmff = nl_shr_mem_2_acc_1_rmff[1:0];
  assign shr_mem_2_cns_PC1 = shr_mem_2_cns_S1 & din_2_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_2_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_2_cns_douta_sho0,
      shr_mem_2_cns_douta_sho1, shr_mem_2_cns_ppidx);
  assign din_2_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_2_cns_douta_sho0,
      shr_mem_2_cns_douta_sho1, shr_mem_2_cns_ppidx_1);
  assign shr_mem_2_cns_addra_shi0 = shr_mem_2_shr_mem_2_mux_3_cse_pff;
  assign shr_mem_2_cns_S1 = (shr_mem_2_cns_ppown_1!=2'b00);
  assign shr_mem_2_cns_S1_pff = (shr_mem_2_acc_1_rmff!=2'b00);
  assign shr_mem_2_and_3_cse_pff = shr_mem_2_cns_S1_pff & (~ shr_mem_2_xor_1_rmff);
  assign shr_mem_2_shr_mem_2_mux_3_cse_pff = MUX_v_8_2_2(dout_2_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_2_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_2_and_3_cse_pff);
  assign shr_mem_2_cns_addrb_shi0 = shr_mem_2_shr_mem_2_mux_3_cse_pff;
  assign shr_mem_2_cns_csa_n_shi0 = shr_mem_2_shr_mem_2_or_cse_pff;
  assign din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_2_cns_S0 = ~((shr_mem_2_cns_ppown==2'b10));
  assign shr_mem_2_cns_S0_pff = ~((shr_mem_2_acc_rmff==2'b10));
  assign shr_mem_2_mux_6_nl = MUX_s_1_2_2(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_2_and_3_cse_pff);
  assign shr_mem_2_shr_mem_2_or_cse_pff = (shr_mem_2_mux_6_nl) | (~((shr_mem_2_cns_S0_pff
      & (~ shr_mem_2_xor_rmff)) | shr_mem_2_and_3_cse_pff));
  assign shr_mem_2_cns_csb_n_shi0 = shr_mem_2_shr_mem_2_or_cse_pff;
  assign shr_mem_2_cns_dinb_shi0 = MUX_v_64_2_2(dout_2_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_2_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_2_and_3_cse_pff);
  assign shr_mem_2_cns_addra_shi1 = shr_mem_2_shr_mem_2_mux_2_cse_pff;
  assign shr_mem_2_and_5_cse_pff = shr_mem_2_cns_S1_pff & shr_mem_2_xor_1_rmff;
  assign shr_mem_2_shr_mem_2_mux_2_cse_pff = MUX_v_8_2_2(dout_2_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_2_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_2_and_5_cse_pff);
  assign shr_mem_2_cns_addrb_shi1 = shr_mem_2_shr_mem_2_mux_2_cse_pff;
  assign shr_mem_2_cns_csa_n_shi1 = shr_mem_2_shr_mem_2_or_1_cse_pff;
  assign shr_mem_2_mux_7_nl = MUX_s_1_2_2(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_2_and_5_cse_pff);
  assign shr_mem_2_shr_mem_2_or_1_cse_pff = (shr_mem_2_mux_7_nl) | (~((shr_mem_2_cns_S0_pff
      & shr_mem_2_xor_rmff) | shr_mem_2_and_5_cse_pff));
  assign shr_mem_2_cns_csb_n_shi1 = shr_mem_2_shr_mem_2_or_1_cse_pff;
  assign shr_mem_2_cns_dinb_shi1 = MUX_v_64_2_2(dout_2_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_2_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_2_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_2_cns_ppidx <= 1'b0;
      shr_mem_2_cns_ppown <= 2'b0;
      shr_mem_2_cns_ppidx_1 <= 1'b0;
      shr_mem_2_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_2_cns_ppidx <= shr_mem_2_xor_rmff;
      shr_mem_2_cns_ppown <= shr_mem_2_acc_rmff;
      shr_mem_2_cns_ppidx_1 <= shr_mem_2_xor_1_rmff;
      shr_mem_2_cns_ppown_1 <= shr_mem_2_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeYeetf_1_cns_bctl
// ------------------------------------------------------------------


module double_buffeYeetf_1_cns_bctl (
  clk, rst, dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_1_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_1_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_1_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_1_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_1_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_1_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_1_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_1_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_1_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_1_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_1_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_1_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_1_cns_S0, shr_mem_1_cns_R0, shr_mem_1_cns_S1, shr_mem_1_cns_R1, shr_mem_1_cns_addra_shi0,
      shr_mem_1_cns_addra_shi1, shr_mem_1_cns_addrb_shi0, shr_mem_1_cns_addrb_shi1,
      shr_mem_1_cns_csa_n_shi0, shr_mem_1_cns_csa_n_shi1, shr_mem_1_cns_csb_n_shi0,
      shr_mem_1_cns_csb_n_shi1, shr_mem_1_cns_dinb_shi0, shr_mem_1_cns_dinb_shi1,
      shr_mem_1_cns_douta_sho0, shr_mem_1_cns_douta_sho1, shr_mem_1_cns_S1_pff, din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff, shr_mem_1_cns_S0_pff
);
  input clk;
  input rst;
  input dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_1_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_1_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_1_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_1_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_1_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_1_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_1_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_1_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_1_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_1_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_1_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  output din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_1_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_1_cns_S0;
  input shr_mem_1_cns_R0;
  output shr_mem_1_cns_S1;
  input shr_mem_1_cns_R1;
  output [7:0] shr_mem_1_cns_addra_shi0;
  output [7:0] shr_mem_1_cns_addra_shi1;
  output [7:0] shr_mem_1_cns_addrb_shi0;
  output [7:0] shr_mem_1_cns_addrb_shi1;
  output shr_mem_1_cns_csa_n_shi0;
  output shr_mem_1_cns_csa_n_shi1;
  output shr_mem_1_cns_csb_n_shi0;
  output shr_mem_1_cns_csb_n_shi1;
  output [63:0] shr_mem_1_cns_dinb_shi0;
  output [63:0] shr_mem_1_cns_dinb_shi1;
  input [63:0] shr_mem_1_cns_douta_sho0;
  input [63:0] shr_mem_1_cns_douta_sho1;
  output shr_mem_1_cns_S1_pff;
  input din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  input dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  output dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output shr_mem_1_cns_S0_pff;


  // Interconnect Declarations
  reg dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  reg din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  wire shr_mem_1_cns_PC0;
  reg shr_mem_1_cns_ppidx;
  reg [1:0] shr_mem_1_cns_ppown;
  wire shr_mem_1_cns_PC1;
  reg shr_mem_1_cns_ppidx_1;
  reg [1:0] shr_mem_1_cns_ppown_1;
  wire [7:0] shr_mem_1_shr_mem_1_mux_3_cse_pff;
  wire shr_mem_1_and_3_cse_pff;
  wire [1:0] shr_mem_1_acc_1_rmff;
  wire [3:0] nl_shr_mem_1_acc_1_rmff;
  wire shr_mem_1_xor_1_rmff;
  wire shr_mem_1_shr_mem_1_or_cse_pff;
  wire [1:0] shr_mem_1_acc_rmff;
  wire [3:0] nl_shr_mem_1_acc_rmff;
  wire shr_mem_1_xor_rmff;
  wire [7:0] shr_mem_1_shr_mem_1_mux_2_cse_pff;
  wire shr_mem_1_and_5_cse_pff;
  wire shr_mem_1_shr_mem_1_or_1_cse_pff;

  wire[0:0] shr_mem_1_mux_6_nl;
  wire[0:0] shr_mem_1_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_1_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_1_cns_R0;
  assign din_1_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_1_cns_R1;
  assign shr_mem_1_xor_rmff = shr_mem_1_cns_ppidx ^ shr_mem_1_cns_PC0;
  assign nl_shr_mem_1_acc_rmff = shr_mem_1_cns_ppown + conv_u2u_1_2(shr_mem_1_cns_PC0)
      + conv_s2u_1_2(shr_mem_1_cns_PC1);
  assign shr_mem_1_acc_rmff = nl_shr_mem_1_acc_rmff[1:0];
  assign shr_mem_1_cns_PC0 = shr_mem_1_cns_S0 & dout_1_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_1_xor_1_rmff = shr_mem_1_cns_ppidx_1 ^ shr_mem_1_cns_PC1;
  assign nl_shr_mem_1_acc_1_rmff = shr_mem_1_cns_ppown_1 + conv_u2u_1_2(shr_mem_1_cns_PC1)
      + conv_s2u_1_2(shr_mem_1_cns_PC0);
  assign shr_mem_1_acc_1_rmff = nl_shr_mem_1_acc_1_rmff[1:0];
  assign shr_mem_1_cns_PC1 = shr_mem_1_cns_S1 & din_1_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_1_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_1_cns_douta_sho0,
      shr_mem_1_cns_douta_sho1, shr_mem_1_cns_ppidx);
  assign din_1_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_1_cns_douta_sho0,
      shr_mem_1_cns_douta_sho1, shr_mem_1_cns_ppidx_1);
  assign shr_mem_1_cns_addra_shi0 = shr_mem_1_shr_mem_1_mux_3_cse_pff;
  assign shr_mem_1_cns_S1 = (shr_mem_1_cns_ppown_1!=2'b00);
  assign shr_mem_1_cns_S1_pff = (shr_mem_1_acc_1_rmff!=2'b00);
  assign shr_mem_1_and_3_cse_pff = shr_mem_1_cns_S1_pff & (~ shr_mem_1_xor_1_rmff);
  assign shr_mem_1_shr_mem_1_mux_3_cse_pff = MUX_v_8_2_2(dout_1_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_1_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_1_and_3_cse_pff);
  assign shr_mem_1_cns_addrb_shi0 = shr_mem_1_shr_mem_1_mux_3_cse_pff;
  assign shr_mem_1_cns_csa_n_shi0 = shr_mem_1_shr_mem_1_or_cse_pff;
  assign din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff = din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud = ~ dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy;
  assign dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff =
      dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign shr_mem_1_cns_S0 = ~((shr_mem_1_cns_ppown==2'b10));
  assign shr_mem_1_cns_S0_pff = ~((shr_mem_1_acc_rmff==2'b10));
  assign shr_mem_1_mux_6_nl = MUX_s_1_2_2(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_1_and_3_cse_pff);
  assign shr_mem_1_shr_mem_1_or_cse_pff = (shr_mem_1_mux_6_nl) | (~((shr_mem_1_cns_S0_pff
      & (~ shr_mem_1_xor_rmff)) | shr_mem_1_and_3_cse_pff));
  assign shr_mem_1_cns_csb_n_shi0 = shr_mem_1_shr_mem_1_or_cse_pff;
  assign shr_mem_1_cns_dinb_shi0 = MUX_v_64_2_2(dout_1_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_1_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_1_and_3_cse_pff);
  assign shr_mem_1_cns_addra_shi1 = shr_mem_1_shr_mem_1_mux_2_cse_pff;
  assign shr_mem_1_and_5_cse_pff = shr_mem_1_cns_S1_pff & shr_mem_1_xor_1_rmff;
  assign shr_mem_1_shr_mem_1_mux_2_cse_pff = MUX_v_8_2_2(dout_1_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_1_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_1_and_5_cse_pff);
  assign shr_mem_1_cns_addrb_shi1 = shr_mem_1_shr_mem_1_mux_2_cse_pff;
  assign shr_mem_1_cns_csa_n_shi1 = shr_mem_1_shr_mem_1_or_1_cse_pff;
  assign shr_mem_1_mux_7_nl = MUX_s_1_2_2(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff,
      din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, shr_mem_1_and_5_cse_pff);
  assign shr_mem_1_shr_mem_1_or_1_cse_pff = (shr_mem_1_mux_7_nl) | (~((shr_mem_1_cns_S0_pff
      & shr_mem_1_xor_rmff) | shr_mem_1_and_5_cse_pff));
  assign shr_mem_1_cns_csb_n_shi1 = shr_mem_1_shr_mem_1_or_1_cse_pff;
  assign shr_mem_1_cns_dinb_shi1 = MUX_v_64_2_2(dout_1_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_1_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_1_and_5_cse_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= 1'b0;
      shr_mem_1_cns_ppidx <= 1'b0;
      shr_mem_1_cns_ppown <= 2'b0;
      shr_mem_1_cns_ppidx_1 <= 1'b0;
      shr_mem_1_cns_ppown_1 <= 2'b0;
    end
    else begin
      dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buy <= ~ din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
      shr_mem_1_cns_ppidx <= shr_mem_1_xor_rmff;
      shr_mem_1_cns_ppown <= shr_mem_1_acc_rmff;
      shr_mem_1_cns_ppidx_1 <= shr_mem_1_xor_1_rmff;
      shr_mem_1_cns_ppown_1 <= shr_mem_1_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffeYeetf_0_cns_bctl
// ------------------------------------------------------------------


module double_buffeYeetf_0_cns_bctl (
  clk, rst, din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_0_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_0_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_0_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_0_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_0_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_0_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, dout_0_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, din_0_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_0_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_0_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_0_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_0_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_0_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_0_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz, din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz,
      din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_0_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_0_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_1_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_1_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_2_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_2_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_3_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_3_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_4_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_4_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_5_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_5_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_6_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_6_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_7_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_7_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_8_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_8_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_9_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_9_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_10_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_10_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_11_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_11_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_12_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_12_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_13_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_13_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_14_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_14_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, dout_15_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud, din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud,
      din_15_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud, dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud,
      shr_mem_0_cns_S0, shr_mem_0_cns_R0, shr_mem_0_cns_S1, shr_mem_0_cns_R1, shr_mem_0_cns_addra_shi0,
      shr_mem_0_cns_addra_shi1, shr_mem_0_cns_addrb_shi0, shr_mem_0_cns_addrb_shi1,
      shr_mem_0_cns_csa_n_shi0, shr_mem_0_cns_csa_n_shi1, shr_mem_0_cns_csb_n_shi0,
      shr_mem_0_cns_csb_n_shi1, shr_mem_0_cns_dinb_shi0, shr_mem_0_cns_dinb_shi1,
      shr_mem_0_cns_douta_sho0, shr_mem_0_cns_douta_sho1, shr_mem_0_cns_S1_pff, shr_mem_0_cns_S0_pff,
      din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff,
      dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff, dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff
);
  input clk;
  input rst;
  output din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_0_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input dout_0_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_0_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] dout_0_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] dout_0_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] dout_0_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_0_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_0_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input din_0_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_0_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [7:0] din_0_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  input [63:0] din_0_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output [63:0] din_0_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_0_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  output din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  output din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  input din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_0_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_0_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_1_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_1_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_2_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_2_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_3_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_3_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_4_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_4_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_5_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_5_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_6_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_6_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_7_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_7_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_8_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_8_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_9_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_9_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_10_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_10_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_11_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_11_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_12_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_12_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_13_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_13_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_14_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_14_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input dout_15_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  input din_15_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  input dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  output shr_mem_0_cns_S0;
  input shr_mem_0_cns_R0;
  output shr_mem_0_cns_S1;
  input shr_mem_0_cns_R1;
  output [7:0] shr_mem_0_cns_addra_shi0;
  output [7:0] shr_mem_0_cns_addra_shi1;
  output [7:0] shr_mem_0_cns_addrb_shi0;
  output [7:0] shr_mem_0_cns_addrb_shi1;
  output shr_mem_0_cns_csa_n_shi0;
  output shr_mem_0_cns_csa_n_shi1;
  output shr_mem_0_cns_csb_n_shi0;
  output shr_mem_0_cns_csb_n_shi1;
  output [63:0] shr_mem_0_cns_dinb_shi0;
  output [63:0] shr_mem_0_cns_dinb_shi1;
  input [63:0] shr_mem_0_cns_douta_sho0;
  input [63:0] shr_mem_0_cns_douta_sho1;
  output shr_mem_0_cns_S1_pff;
  output shr_mem_0_cns_S0_pff;
  output din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  output dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff;
  input dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;


  // Interconnect Declarations
  wire shr_mem_0_cns_PC0;
  reg shr_mem_0_cns_ppidx;
  reg [1:0] shr_mem_0_cns_ppown;
  wire shr_mem_0_cns_PC1;
  reg shr_mem_0_cns_ppidx_1;
  reg [1:0] shr_mem_0_cns_ppown_1;
  wire [7:0] shr_mem_0_shr_mem_0_mux_3_cse_pff;
  wire shr_mem_0_and_3_cse_pff;
  wire [1:0] shr_mem_0_acc_1_rmff;
  wire [3:0] nl_shr_mem_0_acc_1_rmff;
  wire shr_mem_0_xor_1_rmff;
  wire shr_mem_0_shr_mem_0_shr_mem_0_nand_cse_pff;
  wire [1:0] shr_mem_0_acc_rmff;
  wire [3:0] nl_shr_mem_0_acc_rmff;
  wire shr_mem_0_xor_rmff;
  wire [7:0] shr_mem_0_shr_mem_0_mux_2_cse_pff;
  wire shr_mem_0_and_5_cse_pff;
  wire shr_mem_0_shr_mem_0_shr_mem_0_nand_1_cse_pff;

  wire[0:0] shr_mem_0_mux_6_nl;
  wire[0:0] shr_mem_0_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_0_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_0_cns_R0;
  assign din_0_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = shr_mem_0_cns_R1;
  assign shr_mem_0_xor_rmff = shr_mem_0_cns_ppidx ^ shr_mem_0_cns_PC0;
  assign nl_shr_mem_0_acc_rmff = shr_mem_0_cns_ppown + conv_u2u_1_2(shr_mem_0_cns_PC0)
      + conv_s2u_1_2(shr_mem_0_cns_PC1);
  assign shr_mem_0_acc_rmff = nl_shr_mem_0_acc_rmff[1:0];
  assign shr_mem_0_cns_PC0 = shr_mem_0_cns_S0 & dout_0_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign shr_mem_0_xor_1_rmff = shr_mem_0_cns_ppidx_1 ^ shr_mem_0_cns_PC1;
  assign nl_shr_mem_0_acc_1_rmff = shr_mem_0_cns_ppown_1 + conv_u2u_1_2(shr_mem_0_cns_PC1)
      + conv_s2u_1_2(shr_mem_0_cns_PC0);
  assign shr_mem_0_acc_1_rmff = nl_shr_mem_0_acc_1_rmff[1:0];
  assign shr_mem_0_cns_PC1 = shr_mem_0_cns_S1 & din_0_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  assign dout_0_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_0_cns_douta_sho0,
      shr_mem_0_cns_douta_sho1, shr_mem_0_cns_ppidx);
  assign din_0_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst = MUX_v_64_2_2(shr_mem_0_cns_douta_sho0,
      shr_mem_0_cns_douta_sho1, shr_mem_0_cns_ppidx_1);
  assign shr_mem_0_cns_addra_shi0 = shr_mem_0_shr_mem_0_mux_3_cse_pff;
  assign shr_mem_0_cns_S1 = (shr_mem_0_cns_ppown_1!=2'b00);
  assign shr_mem_0_cns_S1_pff = (shr_mem_0_acc_1_rmff!=2'b00);
  assign shr_mem_0_and_3_cse_pff = shr_mem_0_cns_S1_pff & (~ shr_mem_0_xor_1_rmff);
  assign shr_mem_0_shr_mem_0_mux_3_cse_pff = MUX_v_8_2_2(dout_0_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_0_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_0_and_3_cse_pff);
  assign shr_mem_0_cns_addrb_shi0 = shr_mem_0_shr_mem_0_mux_3_cse_pff;
  assign shr_mem_0_cns_csa_n_shi0 = shr_mem_0_shr_mem_0_shr_mem_0_nand_cse_pff;
  assign shr_mem_0_cns_S0 = ~((shr_mem_0_cns_ppown==2'b10));
  assign shr_mem_0_cns_S0_pff = ~((shr_mem_0_acc_rmff==2'b10));
  assign shr_mem_0_mux_6_nl = MUX_s_1_2_2(dout_0_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_0_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_0_and_3_cse_pff);
  assign shr_mem_0_shr_mem_0_shr_mem_0_nand_cse_pff = (shr_mem_0_mux_6_nl) | (~((shr_mem_0_cns_S0_pff
      & (~ shr_mem_0_xor_rmff)) | shr_mem_0_and_3_cse_pff));
  assign shr_mem_0_cns_csb_n_shi0 = shr_mem_0_shr_mem_0_shr_mem_0_nand_cse_pff;
  assign shr_mem_0_cns_dinb_shi0 = MUX_v_64_2_2(dout_0_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_0_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_0_and_3_cse_pff);
  assign shr_mem_0_cns_addra_shi1 = shr_mem_0_shr_mem_0_mux_2_cse_pff;
  assign shr_mem_0_and_5_cse_pff = shr_mem_0_cns_S1_pff & shr_mem_0_xor_1_rmff;
  assign shr_mem_0_shr_mem_0_mux_2_cse_pff = MUX_v_8_2_2(dout_0_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_0_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_0_and_5_cse_pff);
  assign shr_mem_0_cns_addrb_shi1 = shr_mem_0_shr_mem_0_mux_2_cse_pff;
  assign shr_mem_0_cns_csa_n_shi1 = shr_mem_0_shr_mem_0_shr_mem_0_nand_1_cse_pff;
  assign shr_mem_0_mux_7_nl = MUX_s_1_2_2(dout_0_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_0_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_0_and_5_cse_pff);
  assign shr_mem_0_shr_mem_0_shr_mem_0_nand_1_cse_pff = (shr_mem_0_mux_7_nl) | (~((shr_mem_0_cns_S0_pff
      & shr_mem_0_xor_rmff) | shr_mem_0_and_5_cse_pff));
  assign shr_mem_0_cns_csb_n_shi1 = shr_mem_0_shr_mem_0_shr_mem_0_nand_1_cse_pff;
  assign shr_mem_0_cns_dinb_shi1 = MUX_v_64_2_2(dout_0_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst,
      din_0_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst, shr_mem_0_and_5_cse_pff);
  assign din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  assign dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz = dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  assign dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff = dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff;
  always @(posedge clk) begin
    if ( rst ) begin
      shr_mem_0_cns_ppidx <= 1'b0;
      shr_mem_0_cns_ppown <= 2'b0;
      shr_mem_0_cns_ppidx_1 <= 1'b0;
      shr_mem_0_cns_ppown_1 <= 2'b0;
    end
    else begin
      shr_mem_0_cns_ppidx <= shr_mem_0_xor_rmff;
      shr_mem_0_cns_ppown <= shr_mem_0_acc_rmff;
      shr_mem_0_cns_ppidx_1 <= shr_mem_0_xor_1_rmff;
      shr_mem_0_cns_ppown_1 <= shr_mem_0_acc_1_rmff;
    end
  end

  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function  [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function  [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    unreg_hier_31
// ------------------------------------------------------------------


module unreg_hier_31 (
  in_0, out_0
);
  input in_0;
  output out_0;



  // Interconnect Declarations for Component Instantiations 
  assign out_0 = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_128_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_128_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_15_and_nl;
  wire dout_15_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_15_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_15_and_nl);
  assign dout_15_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_15_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_127_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_127_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_14_and_nl;
  wire dout_14_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_14_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_14_and_nl);
  assign dout_14_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_14_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_126_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_126_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_13_and_nl;
  wire dout_13_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_13_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_13_and_nl);
  assign dout_13_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_13_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_125_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_125_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_12_and_nl;
  wire dout_12_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_12_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_12_and_nl);
  assign dout_12_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_12_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_124_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_124_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_11_and_nl;
  wire dout_11_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_11_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_11_and_nl);
  assign dout_11_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_11_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_123_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_123_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_10_and_nl;
  wire dout_10_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_10_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_10_and_nl);
  assign dout_10_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_10_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_122_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_122_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_9_and_nl;
  wire dout_9_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_9_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_9_and_nl);
  assign dout_9_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_9_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_121_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_121_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_8_and_nl;
  wire dout_8_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_8_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_8_and_nl);
  assign dout_8_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_8_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_120_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_120_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_7_and_nl;
  wire dout_7_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_7_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_7_and_nl);
  assign dout_7_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_7_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_119_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_119_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_6_and_nl;
  wire dout_6_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_6_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_6_and_nl);
  assign dout_6_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_6_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_118_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_118_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_5_and_nl;
  wire dout_5_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_5_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_5_and_nl);
  assign dout_5_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_5_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_117_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_117_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_4_and_nl;
  wire dout_4_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_4_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_4_and_nl);
  assign dout_4_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_4_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_116_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_116_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_3_and_nl;
  wire dout_3_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_3_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_3_and_nl);
  assign dout_3_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_3_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_115_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_115_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_2_and_nl;
  wire dout_2_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_2_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_2_and_nl);
  assign dout_2_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_2_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_114_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_114_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_1_and_nl;
  wire dout_1_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_1_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_1_and_nl);
  assign dout_1_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_1_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_113_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_113_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_0_and_nl;
  wire dout_0_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign dout_0_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (dout_0_and_nl);
  assign dout_0_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (dout_0_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_staller
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_staller (
  clk, rst, core_wen, din_rsci_wen_comp, core_wten, dout_15_rsc_req_obj_wen_comp,
      dout_14_rsc_req_obj_wen_comp, dout_13_rsc_req_obj_wen_comp, dout_12_rsc_req_obj_wen_comp,
      dout_11_rsc_req_obj_wen_comp, dout_10_rsc_req_obj_wen_comp, dout_9_rsc_req_obj_wen_comp,
      dout_8_rsc_req_obj_wen_comp, dout_7_rsc_req_obj_wen_comp, dout_6_rsc_req_obj_wen_comp,
      dout_5_rsc_req_obj_wen_comp, dout_4_rsc_req_obj_wen_comp, dout_3_rsc_req_obj_wen_comp,
      dout_2_rsc_req_obj_wen_comp, dout_1_rsc_req_obj_wen_comp, dout_0_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  input din_rsci_wen_comp;
  output core_wten;
  input dout_15_rsc_req_obj_wen_comp;
  input dout_14_rsc_req_obj_wen_comp;
  input dout_13_rsc_req_obj_wen_comp;
  input dout_12_rsc_req_obj_wen_comp;
  input dout_11_rsc_req_obj_wen_comp;
  input dout_10_rsc_req_obj_wen_comp;
  input dout_9_rsc_req_obj_wen_comp;
  input dout_8_rsc_req_obj_wen_comp;
  input dout_7_rsc_req_obj_wen_comp;
  input dout_6_rsc_req_obj_wen_comp;
  input dout_5_rsc_req_obj_wen_comp;
  input dout_4_rsc_req_obj_wen_comp;
  input dout_3_rsc_req_obj_wen_comp;
  input dout_2_rsc_req_obj_wen_comp;
  input dout_1_rsc_req_obj_wen_comp;
  input dout_0_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = din_rsci_wen_comp & dout_15_rsc_req_obj_wen_comp & dout_14_rsc_req_obj_wen_comp
      & dout_13_rsc_req_obj_wen_comp & dout_12_rsc_req_obj_wen_comp & dout_11_rsc_req_obj_wen_comp
      & dout_10_rsc_req_obj_wen_comp & dout_9_rsc_req_obj_wen_comp & dout_8_rsc_req_obj_wen_comp
      & dout_7_rsc_req_obj_wen_comp & dout_6_rsc_req_obj_wen_comp & dout_5_rsc_req_obj_wen_comp
      & dout_4_rsc_req_obj_wen_comp & dout_3_rsc_req_obj_wen_comp & dout_2_rsc_req_obj_wen_comp
      & dout_1_rsc_req_obj_wen_comp & dout_0_rsc_req_obj_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_dp
    (
  clk, rst, dout_0_rsc_req_obj_oswt, dout_0_rsc_req_obj_wen_comp, dout_0_rsc_req_obj_biwt,
      dout_0_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_0_rsc_req_obj_oswt;
  output dout_0_rsc_req_obj_wen_comp;
  input dout_0_rsc_req_obj_biwt;
  input dout_0_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_0_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_0_rsc_req_obj_wen_comp = (~ dout_0_rsc_req_obj_oswt) | dout_0_rsc_req_obj_biwt
      | dout_0_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_0_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_0_rsc_req_obj_bcwt <= ~((~(dout_0_rsc_req_obj_bcwt | dout_0_rsc_req_obj_biwt))
          | dout_0_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_0_rsc_req_obj_oswt, dout_0_rsc_req_obj_vd,
      dout_0_rsc_req_obj_biwt, dout_0_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_0_rsc_req_obj_oswt;
  input dout_0_rsc_req_obj_vd;
  output dout_0_rsc_req_obj_biwt;
  output dout_0_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_0_rsc_req_obj_pdswt0;
  reg dout_0_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_0_rsc_req_obj_pdswt0 = (~ core_wten) & dout_0_rsc_req_obj_oswt;
  assign dout_0_rsc_req_obj_biwt = (dout_0_rsc_req_obj_pdswt0 | dout_0_rsc_req_obj_icwt)
      & dout_0_rsc_req_obj_vd;
  assign dout_0_rsc_req_obj_bdwt = dout_0_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_0_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_0_rsc_req_obj_icwt <= ~((~(dout_0_rsc_req_obj_icwt | dout_0_rsc_req_obj_pdswt0))
          | dout_0_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_dp
    (
  clk, rst, dout_1_rsc_req_obj_oswt, dout_1_rsc_req_obj_wen_comp, dout_1_rsc_req_obj_biwt,
      dout_1_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_1_rsc_req_obj_oswt;
  output dout_1_rsc_req_obj_wen_comp;
  input dout_1_rsc_req_obj_biwt;
  input dout_1_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_1_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_1_rsc_req_obj_wen_comp = (~ dout_1_rsc_req_obj_oswt) | dout_1_rsc_req_obj_biwt
      | dout_1_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_1_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_1_rsc_req_obj_bcwt <= ~((~(dout_1_rsc_req_obj_bcwt | dout_1_rsc_req_obj_biwt))
          | dout_1_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_1_rsc_req_obj_oswt, dout_1_rsc_req_obj_vd,
      dout_1_rsc_req_obj_biwt, dout_1_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_1_rsc_req_obj_oswt;
  input dout_1_rsc_req_obj_vd;
  output dout_1_rsc_req_obj_biwt;
  output dout_1_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_1_rsc_req_obj_pdswt0;
  reg dout_1_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_1_rsc_req_obj_pdswt0 = (~ core_wten) & dout_1_rsc_req_obj_oswt;
  assign dout_1_rsc_req_obj_biwt = (dout_1_rsc_req_obj_pdswt0 | dout_1_rsc_req_obj_icwt)
      & dout_1_rsc_req_obj_vd;
  assign dout_1_rsc_req_obj_bdwt = dout_1_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_1_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_1_rsc_req_obj_icwt <= ~((~(dout_1_rsc_req_obj_icwt | dout_1_rsc_req_obj_pdswt0))
          | dout_1_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_dp
    (
  clk, rst, dout_2_rsc_req_obj_oswt, dout_2_rsc_req_obj_wen_comp, dout_2_rsc_req_obj_biwt,
      dout_2_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_2_rsc_req_obj_oswt;
  output dout_2_rsc_req_obj_wen_comp;
  input dout_2_rsc_req_obj_biwt;
  input dout_2_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_2_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_2_rsc_req_obj_wen_comp = (~ dout_2_rsc_req_obj_oswt) | dout_2_rsc_req_obj_biwt
      | dout_2_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_2_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_2_rsc_req_obj_bcwt <= ~((~(dout_2_rsc_req_obj_bcwt | dout_2_rsc_req_obj_biwt))
          | dout_2_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_2_rsc_req_obj_oswt, dout_2_rsc_req_obj_vd,
      dout_2_rsc_req_obj_biwt, dout_2_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_2_rsc_req_obj_oswt;
  input dout_2_rsc_req_obj_vd;
  output dout_2_rsc_req_obj_biwt;
  output dout_2_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_2_rsc_req_obj_pdswt0;
  reg dout_2_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_2_rsc_req_obj_pdswt0 = (~ core_wten) & dout_2_rsc_req_obj_oswt;
  assign dout_2_rsc_req_obj_biwt = (dout_2_rsc_req_obj_pdswt0 | dout_2_rsc_req_obj_icwt)
      & dout_2_rsc_req_obj_vd;
  assign dout_2_rsc_req_obj_bdwt = dout_2_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_2_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_2_rsc_req_obj_icwt <= ~((~(dout_2_rsc_req_obj_icwt | dout_2_rsc_req_obj_pdswt0))
          | dout_2_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_dp
    (
  clk, rst, dout_3_rsc_req_obj_oswt, dout_3_rsc_req_obj_wen_comp, dout_3_rsc_req_obj_biwt,
      dout_3_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_3_rsc_req_obj_oswt;
  output dout_3_rsc_req_obj_wen_comp;
  input dout_3_rsc_req_obj_biwt;
  input dout_3_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_3_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_3_rsc_req_obj_wen_comp = (~ dout_3_rsc_req_obj_oswt) | dout_3_rsc_req_obj_biwt
      | dout_3_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_3_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_3_rsc_req_obj_bcwt <= ~((~(dout_3_rsc_req_obj_bcwt | dout_3_rsc_req_obj_biwt))
          | dout_3_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_3_rsc_req_obj_oswt, dout_3_rsc_req_obj_vd,
      dout_3_rsc_req_obj_biwt, dout_3_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_3_rsc_req_obj_oswt;
  input dout_3_rsc_req_obj_vd;
  output dout_3_rsc_req_obj_biwt;
  output dout_3_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_3_rsc_req_obj_pdswt0;
  reg dout_3_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_3_rsc_req_obj_pdswt0 = (~ core_wten) & dout_3_rsc_req_obj_oswt;
  assign dout_3_rsc_req_obj_biwt = (dout_3_rsc_req_obj_pdswt0 | dout_3_rsc_req_obj_icwt)
      & dout_3_rsc_req_obj_vd;
  assign dout_3_rsc_req_obj_bdwt = dout_3_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_3_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_3_rsc_req_obj_icwt <= ~((~(dout_3_rsc_req_obj_icwt | dout_3_rsc_req_obj_pdswt0))
          | dout_3_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_dp
    (
  clk, rst, dout_4_rsc_req_obj_oswt, dout_4_rsc_req_obj_wen_comp, dout_4_rsc_req_obj_biwt,
      dout_4_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_4_rsc_req_obj_oswt;
  output dout_4_rsc_req_obj_wen_comp;
  input dout_4_rsc_req_obj_biwt;
  input dout_4_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_4_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_4_rsc_req_obj_wen_comp = (~ dout_4_rsc_req_obj_oswt) | dout_4_rsc_req_obj_biwt
      | dout_4_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_4_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_4_rsc_req_obj_bcwt <= ~((~(dout_4_rsc_req_obj_bcwt | dout_4_rsc_req_obj_biwt))
          | dout_4_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_4_rsc_req_obj_oswt, dout_4_rsc_req_obj_vd,
      dout_4_rsc_req_obj_biwt, dout_4_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_4_rsc_req_obj_oswt;
  input dout_4_rsc_req_obj_vd;
  output dout_4_rsc_req_obj_biwt;
  output dout_4_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_4_rsc_req_obj_pdswt0;
  reg dout_4_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_4_rsc_req_obj_pdswt0 = (~ core_wten) & dout_4_rsc_req_obj_oswt;
  assign dout_4_rsc_req_obj_biwt = (dout_4_rsc_req_obj_pdswt0 | dout_4_rsc_req_obj_icwt)
      & dout_4_rsc_req_obj_vd;
  assign dout_4_rsc_req_obj_bdwt = dout_4_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_4_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_4_rsc_req_obj_icwt <= ~((~(dout_4_rsc_req_obj_icwt | dout_4_rsc_req_obj_pdswt0))
          | dout_4_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_dp
    (
  clk, rst, dout_5_rsc_req_obj_oswt, dout_5_rsc_req_obj_wen_comp, dout_5_rsc_req_obj_biwt,
      dout_5_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_5_rsc_req_obj_oswt;
  output dout_5_rsc_req_obj_wen_comp;
  input dout_5_rsc_req_obj_biwt;
  input dout_5_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_5_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_5_rsc_req_obj_wen_comp = (~ dout_5_rsc_req_obj_oswt) | dout_5_rsc_req_obj_biwt
      | dout_5_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_5_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_5_rsc_req_obj_bcwt <= ~((~(dout_5_rsc_req_obj_bcwt | dout_5_rsc_req_obj_biwt))
          | dout_5_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_5_rsc_req_obj_oswt, dout_5_rsc_req_obj_vd,
      dout_5_rsc_req_obj_biwt, dout_5_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_5_rsc_req_obj_oswt;
  input dout_5_rsc_req_obj_vd;
  output dout_5_rsc_req_obj_biwt;
  output dout_5_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_5_rsc_req_obj_pdswt0;
  reg dout_5_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_5_rsc_req_obj_pdswt0 = (~ core_wten) & dout_5_rsc_req_obj_oswt;
  assign dout_5_rsc_req_obj_biwt = (dout_5_rsc_req_obj_pdswt0 | dout_5_rsc_req_obj_icwt)
      & dout_5_rsc_req_obj_vd;
  assign dout_5_rsc_req_obj_bdwt = dout_5_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_5_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_5_rsc_req_obj_icwt <= ~((~(dout_5_rsc_req_obj_icwt | dout_5_rsc_req_obj_pdswt0))
          | dout_5_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_dp
    (
  clk, rst, dout_6_rsc_req_obj_oswt, dout_6_rsc_req_obj_wen_comp, dout_6_rsc_req_obj_biwt,
      dout_6_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_6_rsc_req_obj_oswt;
  output dout_6_rsc_req_obj_wen_comp;
  input dout_6_rsc_req_obj_biwt;
  input dout_6_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_6_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_6_rsc_req_obj_wen_comp = (~ dout_6_rsc_req_obj_oswt) | dout_6_rsc_req_obj_biwt
      | dout_6_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_6_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_6_rsc_req_obj_bcwt <= ~((~(dout_6_rsc_req_obj_bcwt | dout_6_rsc_req_obj_biwt))
          | dout_6_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_6_rsc_req_obj_oswt, dout_6_rsc_req_obj_vd,
      dout_6_rsc_req_obj_biwt, dout_6_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_6_rsc_req_obj_oswt;
  input dout_6_rsc_req_obj_vd;
  output dout_6_rsc_req_obj_biwt;
  output dout_6_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_6_rsc_req_obj_pdswt0;
  reg dout_6_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_6_rsc_req_obj_pdswt0 = (~ core_wten) & dout_6_rsc_req_obj_oswt;
  assign dout_6_rsc_req_obj_biwt = (dout_6_rsc_req_obj_pdswt0 | dout_6_rsc_req_obj_icwt)
      & dout_6_rsc_req_obj_vd;
  assign dout_6_rsc_req_obj_bdwt = dout_6_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_6_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_6_rsc_req_obj_icwt <= ~((~(dout_6_rsc_req_obj_icwt | dout_6_rsc_req_obj_pdswt0))
          | dout_6_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_dp
    (
  clk, rst, dout_7_rsc_req_obj_oswt, dout_7_rsc_req_obj_wen_comp, dout_7_rsc_req_obj_biwt,
      dout_7_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_7_rsc_req_obj_oswt;
  output dout_7_rsc_req_obj_wen_comp;
  input dout_7_rsc_req_obj_biwt;
  input dout_7_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_7_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_7_rsc_req_obj_wen_comp = (~ dout_7_rsc_req_obj_oswt) | dout_7_rsc_req_obj_biwt
      | dout_7_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_7_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_7_rsc_req_obj_bcwt <= ~((~(dout_7_rsc_req_obj_bcwt | dout_7_rsc_req_obj_biwt))
          | dout_7_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_7_rsc_req_obj_oswt, dout_7_rsc_req_obj_vd,
      dout_7_rsc_req_obj_biwt, dout_7_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_7_rsc_req_obj_oswt;
  input dout_7_rsc_req_obj_vd;
  output dout_7_rsc_req_obj_biwt;
  output dout_7_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_7_rsc_req_obj_pdswt0;
  reg dout_7_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_7_rsc_req_obj_pdswt0 = (~ core_wten) & dout_7_rsc_req_obj_oswt;
  assign dout_7_rsc_req_obj_biwt = (dout_7_rsc_req_obj_pdswt0 | dout_7_rsc_req_obj_icwt)
      & dout_7_rsc_req_obj_vd;
  assign dout_7_rsc_req_obj_bdwt = dout_7_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_7_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_7_rsc_req_obj_icwt <= ~((~(dout_7_rsc_req_obj_icwt | dout_7_rsc_req_obj_pdswt0))
          | dout_7_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_dp
    (
  clk, rst, dout_8_rsc_req_obj_oswt, dout_8_rsc_req_obj_wen_comp, dout_8_rsc_req_obj_biwt,
      dout_8_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_8_rsc_req_obj_oswt;
  output dout_8_rsc_req_obj_wen_comp;
  input dout_8_rsc_req_obj_biwt;
  input dout_8_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_8_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_8_rsc_req_obj_wen_comp = (~ dout_8_rsc_req_obj_oswt) | dout_8_rsc_req_obj_biwt
      | dout_8_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_8_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_8_rsc_req_obj_bcwt <= ~((~(dout_8_rsc_req_obj_bcwt | dout_8_rsc_req_obj_biwt))
          | dout_8_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_8_rsc_req_obj_oswt, dout_8_rsc_req_obj_vd,
      dout_8_rsc_req_obj_biwt, dout_8_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_8_rsc_req_obj_oswt;
  input dout_8_rsc_req_obj_vd;
  output dout_8_rsc_req_obj_biwt;
  output dout_8_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_8_rsc_req_obj_pdswt0;
  reg dout_8_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_8_rsc_req_obj_pdswt0 = (~ core_wten) & dout_8_rsc_req_obj_oswt;
  assign dout_8_rsc_req_obj_biwt = (dout_8_rsc_req_obj_pdswt0 | dout_8_rsc_req_obj_icwt)
      & dout_8_rsc_req_obj_vd;
  assign dout_8_rsc_req_obj_bdwt = dout_8_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_8_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_8_rsc_req_obj_icwt <= ~((~(dout_8_rsc_req_obj_icwt | dout_8_rsc_req_obj_pdswt0))
          | dout_8_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_dp
    (
  clk, rst, dout_9_rsc_req_obj_oswt, dout_9_rsc_req_obj_wen_comp, dout_9_rsc_req_obj_biwt,
      dout_9_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_9_rsc_req_obj_oswt;
  output dout_9_rsc_req_obj_wen_comp;
  input dout_9_rsc_req_obj_biwt;
  input dout_9_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_9_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_9_rsc_req_obj_wen_comp = (~ dout_9_rsc_req_obj_oswt) | dout_9_rsc_req_obj_biwt
      | dout_9_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_9_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_9_rsc_req_obj_bcwt <= ~((~(dout_9_rsc_req_obj_bcwt | dout_9_rsc_req_obj_biwt))
          | dout_9_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_9_rsc_req_obj_oswt, dout_9_rsc_req_obj_vd,
      dout_9_rsc_req_obj_biwt, dout_9_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_9_rsc_req_obj_oswt;
  input dout_9_rsc_req_obj_vd;
  output dout_9_rsc_req_obj_biwt;
  output dout_9_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_9_rsc_req_obj_pdswt0;
  reg dout_9_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_9_rsc_req_obj_pdswt0 = (~ core_wten) & dout_9_rsc_req_obj_oswt;
  assign dout_9_rsc_req_obj_biwt = (dout_9_rsc_req_obj_pdswt0 | dout_9_rsc_req_obj_icwt)
      & dout_9_rsc_req_obj_vd;
  assign dout_9_rsc_req_obj_bdwt = dout_9_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_9_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_9_rsc_req_obj_icwt <= ~((~(dout_9_rsc_req_obj_icwt | dout_9_rsc_req_obj_pdswt0))
          | dout_9_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_dp
    (
  clk, rst, dout_10_rsc_req_obj_oswt, dout_10_rsc_req_obj_wen_comp, dout_10_rsc_req_obj_biwt,
      dout_10_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_10_rsc_req_obj_oswt;
  output dout_10_rsc_req_obj_wen_comp;
  input dout_10_rsc_req_obj_biwt;
  input dout_10_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_10_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_10_rsc_req_obj_wen_comp = (~ dout_10_rsc_req_obj_oswt) | dout_10_rsc_req_obj_biwt
      | dout_10_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_10_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_10_rsc_req_obj_bcwt <= ~((~(dout_10_rsc_req_obj_bcwt | dout_10_rsc_req_obj_biwt))
          | dout_10_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_10_rsc_req_obj_oswt, dout_10_rsc_req_obj_vd,
      dout_10_rsc_req_obj_biwt, dout_10_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_10_rsc_req_obj_oswt;
  input dout_10_rsc_req_obj_vd;
  output dout_10_rsc_req_obj_biwt;
  output dout_10_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_10_rsc_req_obj_pdswt0;
  reg dout_10_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_10_rsc_req_obj_pdswt0 = (~ core_wten) & dout_10_rsc_req_obj_oswt;
  assign dout_10_rsc_req_obj_biwt = (dout_10_rsc_req_obj_pdswt0 | dout_10_rsc_req_obj_icwt)
      & dout_10_rsc_req_obj_vd;
  assign dout_10_rsc_req_obj_bdwt = dout_10_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_10_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_10_rsc_req_obj_icwt <= ~((~(dout_10_rsc_req_obj_icwt | dout_10_rsc_req_obj_pdswt0))
          | dout_10_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_dp
    (
  clk, rst, dout_11_rsc_req_obj_oswt, dout_11_rsc_req_obj_wen_comp, dout_11_rsc_req_obj_biwt,
      dout_11_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_11_rsc_req_obj_oswt;
  output dout_11_rsc_req_obj_wen_comp;
  input dout_11_rsc_req_obj_biwt;
  input dout_11_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_11_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_11_rsc_req_obj_wen_comp = (~ dout_11_rsc_req_obj_oswt) | dout_11_rsc_req_obj_biwt
      | dout_11_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_11_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_11_rsc_req_obj_bcwt <= ~((~(dout_11_rsc_req_obj_bcwt | dout_11_rsc_req_obj_biwt))
          | dout_11_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_11_rsc_req_obj_oswt, dout_11_rsc_req_obj_vd,
      dout_11_rsc_req_obj_biwt, dout_11_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_11_rsc_req_obj_oswt;
  input dout_11_rsc_req_obj_vd;
  output dout_11_rsc_req_obj_biwt;
  output dout_11_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_11_rsc_req_obj_pdswt0;
  reg dout_11_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_11_rsc_req_obj_pdswt0 = (~ core_wten) & dout_11_rsc_req_obj_oswt;
  assign dout_11_rsc_req_obj_biwt = (dout_11_rsc_req_obj_pdswt0 | dout_11_rsc_req_obj_icwt)
      & dout_11_rsc_req_obj_vd;
  assign dout_11_rsc_req_obj_bdwt = dout_11_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_11_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_11_rsc_req_obj_icwt <= ~((~(dout_11_rsc_req_obj_icwt | dout_11_rsc_req_obj_pdswt0))
          | dout_11_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_dp
    (
  clk, rst, dout_12_rsc_req_obj_oswt, dout_12_rsc_req_obj_wen_comp, dout_12_rsc_req_obj_biwt,
      dout_12_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_12_rsc_req_obj_oswt;
  output dout_12_rsc_req_obj_wen_comp;
  input dout_12_rsc_req_obj_biwt;
  input dout_12_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_12_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_12_rsc_req_obj_wen_comp = (~ dout_12_rsc_req_obj_oswt) | dout_12_rsc_req_obj_biwt
      | dout_12_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_12_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_12_rsc_req_obj_bcwt <= ~((~(dout_12_rsc_req_obj_bcwt | dout_12_rsc_req_obj_biwt))
          | dout_12_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_12_rsc_req_obj_oswt, dout_12_rsc_req_obj_vd,
      dout_12_rsc_req_obj_biwt, dout_12_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_12_rsc_req_obj_oswt;
  input dout_12_rsc_req_obj_vd;
  output dout_12_rsc_req_obj_biwt;
  output dout_12_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_12_rsc_req_obj_pdswt0;
  reg dout_12_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_12_rsc_req_obj_pdswt0 = (~ core_wten) & dout_12_rsc_req_obj_oswt;
  assign dout_12_rsc_req_obj_biwt = (dout_12_rsc_req_obj_pdswt0 | dout_12_rsc_req_obj_icwt)
      & dout_12_rsc_req_obj_vd;
  assign dout_12_rsc_req_obj_bdwt = dout_12_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_12_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_12_rsc_req_obj_icwt <= ~((~(dout_12_rsc_req_obj_icwt | dout_12_rsc_req_obj_pdswt0))
          | dout_12_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_dp
    (
  clk, rst, dout_13_rsc_req_obj_oswt, dout_13_rsc_req_obj_wen_comp, dout_13_rsc_req_obj_biwt,
      dout_13_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_13_rsc_req_obj_oswt;
  output dout_13_rsc_req_obj_wen_comp;
  input dout_13_rsc_req_obj_biwt;
  input dout_13_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_13_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_13_rsc_req_obj_wen_comp = (~ dout_13_rsc_req_obj_oswt) | dout_13_rsc_req_obj_biwt
      | dout_13_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_13_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_13_rsc_req_obj_bcwt <= ~((~(dout_13_rsc_req_obj_bcwt | dout_13_rsc_req_obj_biwt))
          | dout_13_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_13_rsc_req_obj_oswt, dout_13_rsc_req_obj_vd,
      dout_13_rsc_req_obj_biwt, dout_13_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_13_rsc_req_obj_oswt;
  input dout_13_rsc_req_obj_vd;
  output dout_13_rsc_req_obj_biwt;
  output dout_13_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_13_rsc_req_obj_pdswt0;
  reg dout_13_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_13_rsc_req_obj_pdswt0 = (~ core_wten) & dout_13_rsc_req_obj_oswt;
  assign dout_13_rsc_req_obj_biwt = (dout_13_rsc_req_obj_pdswt0 | dout_13_rsc_req_obj_icwt)
      & dout_13_rsc_req_obj_vd;
  assign dout_13_rsc_req_obj_bdwt = dout_13_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_13_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_13_rsc_req_obj_icwt <= ~((~(dout_13_rsc_req_obj_icwt | dout_13_rsc_req_obj_pdswt0))
          | dout_13_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_dp
    (
  clk, rst, dout_14_rsc_req_obj_oswt, dout_14_rsc_req_obj_wen_comp, dout_14_rsc_req_obj_biwt,
      dout_14_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_14_rsc_req_obj_oswt;
  output dout_14_rsc_req_obj_wen_comp;
  input dout_14_rsc_req_obj_biwt;
  input dout_14_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_14_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_14_rsc_req_obj_wen_comp = (~ dout_14_rsc_req_obj_oswt) | dout_14_rsc_req_obj_biwt
      | dout_14_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_14_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_14_rsc_req_obj_bcwt <= ~((~(dout_14_rsc_req_obj_bcwt | dout_14_rsc_req_obj_biwt))
          | dout_14_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_14_rsc_req_obj_oswt, dout_14_rsc_req_obj_vd,
      dout_14_rsc_req_obj_biwt, dout_14_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_14_rsc_req_obj_oswt;
  input dout_14_rsc_req_obj_vd;
  output dout_14_rsc_req_obj_biwt;
  output dout_14_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_14_rsc_req_obj_pdswt0;
  reg dout_14_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_14_rsc_req_obj_pdswt0 = (~ core_wten) & dout_14_rsc_req_obj_oswt;
  assign dout_14_rsc_req_obj_biwt = (dout_14_rsc_req_obj_pdswt0 | dout_14_rsc_req_obj_icwt)
      & dout_14_rsc_req_obj_vd;
  assign dout_14_rsc_req_obj_bdwt = dout_14_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_14_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_14_rsc_req_obj_icwt <= ~((~(dout_14_rsc_req_obj_icwt | dout_14_rsc_req_obj_pdswt0))
          | dout_14_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_dp
    (
  clk, rst, dout_15_rsc_req_obj_oswt, dout_15_rsc_req_obj_wen_comp, dout_15_rsc_req_obj_biwt,
      dout_15_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input dout_15_rsc_req_obj_oswt;
  output dout_15_rsc_req_obj_wen_comp;
  input dout_15_rsc_req_obj_biwt;
  input dout_15_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg dout_15_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_15_rsc_req_obj_wen_comp = (~ dout_15_rsc_req_obj_oswt) | dout_15_rsc_req_obj_biwt
      | dout_15_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_15_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_15_rsc_req_obj_bcwt <= ~((~(dout_15_rsc_req_obj_bcwt | dout_15_rsc_req_obj_biwt))
          | dout_15_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, dout_15_rsc_req_obj_oswt, dout_15_rsc_req_obj_vd,
      dout_15_rsc_req_obj_biwt, dout_15_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_15_rsc_req_obj_oswt;
  input dout_15_rsc_req_obj_vd;
  output dout_15_rsc_req_obj_biwt;
  output dout_15_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire dout_15_rsc_req_obj_pdswt0;
  reg dout_15_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_15_rsc_req_obj_pdswt0 = (~ core_wten) & dout_15_rsc_req_obj_oswt;
  assign dout_15_rsc_req_obj_biwt = (dout_15_rsc_req_obj_pdswt0 | dout_15_rsc_req_obj_icwt)
      & dout_15_rsc_req_obj_vd;
  assign dout_15_rsc_req_obj_bdwt = dout_15_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_15_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      dout_15_rsc_req_obj_icwt <= ~((~(dout_15_rsc_req_obj_icwt | dout_15_rsc_req_obj_pdswt0))
          | dout_15_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_rls_obj_dout_0_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_rls_obj_dout_0_rsc_rls_wait_ctrl
    (
  core_wten, dout_0_rsc_rls_obj_iswt0, dout_0_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_0_rsc_rls_obj_iswt0;
  output dout_0_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_0_rsc_rls_obj_ld_core_sct = dout_0_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_rls_obj_dout_1_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_rls_obj_dout_1_rsc_rls_wait_ctrl
    (
  core_wten, dout_1_rsc_rls_obj_iswt0, dout_1_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_1_rsc_rls_obj_iswt0;
  output dout_1_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_1_rsc_rls_obj_ld_core_sct = dout_1_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_rls_obj_dout_2_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_rls_obj_dout_2_rsc_rls_wait_ctrl
    (
  core_wten, dout_2_rsc_rls_obj_iswt0, dout_2_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_2_rsc_rls_obj_iswt0;
  output dout_2_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_2_rsc_rls_obj_ld_core_sct = dout_2_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_rls_obj_dout_3_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_rls_obj_dout_3_rsc_rls_wait_ctrl
    (
  core_wten, dout_3_rsc_rls_obj_iswt0, dout_3_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_3_rsc_rls_obj_iswt0;
  output dout_3_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_3_rsc_rls_obj_ld_core_sct = dout_3_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_rls_obj_dout_4_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_rls_obj_dout_4_rsc_rls_wait_ctrl
    (
  core_wten, dout_4_rsc_rls_obj_iswt0, dout_4_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_4_rsc_rls_obj_iswt0;
  output dout_4_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_4_rsc_rls_obj_ld_core_sct = dout_4_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_rls_obj_dout_5_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_rls_obj_dout_5_rsc_rls_wait_ctrl
    (
  core_wten, dout_5_rsc_rls_obj_iswt0, dout_5_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_5_rsc_rls_obj_iswt0;
  output dout_5_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_5_rsc_rls_obj_ld_core_sct = dout_5_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_rls_obj_dout_6_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_rls_obj_dout_6_rsc_rls_wait_ctrl
    (
  core_wten, dout_6_rsc_rls_obj_iswt0, dout_6_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_6_rsc_rls_obj_iswt0;
  output dout_6_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_6_rsc_rls_obj_ld_core_sct = dout_6_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_rls_obj_dout_7_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_rls_obj_dout_7_rsc_rls_wait_ctrl
    (
  core_wten, dout_7_rsc_rls_obj_iswt0, dout_7_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_7_rsc_rls_obj_iswt0;
  output dout_7_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_7_rsc_rls_obj_ld_core_sct = dout_7_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_rls_obj_dout_8_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_rls_obj_dout_8_rsc_rls_wait_ctrl
    (
  core_wten, dout_8_rsc_rls_obj_iswt0, dout_8_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_8_rsc_rls_obj_iswt0;
  output dout_8_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_8_rsc_rls_obj_ld_core_sct = dout_8_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_rls_obj_dout_9_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_rls_obj_dout_9_rsc_rls_wait_ctrl
    (
  core_wten, dout_9_rsc_rls_obj_iswt0, dout_9_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_9_rsc_rls_obj_iswt0;
  output dout_9_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_9_rsc_rls_obj_ld_core_sct = dout_9_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_rls_obj_dout_10_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_rls_obj_dout_10_rsc_rls_wait_ctrl
    (
  core_wten, dout_10_rsc_rls_obj_iswt0, dout_10_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_10_rsc_rls_obj_iswt0;
  output dout_10_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_10_rsc_rls_obj_ld_core_sct = dout_10_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_rls_obj_dout_11_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_rls_obj_dout_11_rsc_rls_wait_ctrl
    (
  core_wten, dout_11_rsc_rls_obj_iswt0, dout_11_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_11_rsc_rls_obj_iswt0;
  output dout_11_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_11_rsc_rls_obj_ld_core_sct = dout_11_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_rls_obj_dout_12_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_rls_obj_dout_12_rsc_rls_wait_ctrl
    (
  core_wten, dout_12_rsc_rls_obj_iswt0, dout_12_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_12_rsc_rls_obj_iswt0;
  output dout_12_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_12_rsc_rls_obj_ld_core_sct = dout_12_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_rls_obj_dout_13_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_rls_obj_dout_13_rsc_rls_wait_ctrl
    (
  core_wten, dout_13_rsc_rls_obj_iswt0, dout_13_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_13_rsc_rls_obj_iswt0;
  output dout_13_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_13_rsc_rls_obj_ld_core_sct = dout_13_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_rls_obj_dout_14_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_rls_obj_dout_14_rsc_rls_wait_ctrl
    (
  core_wten, dout_14_rsc_rls_obj_iswt0, dout_14_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_14_rsc_rls_obj_iswt0;
  output dout_14_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_14_rsc_rls_obj_ld_core_sct = dout_14_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_rls_obj_dout_15_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_rls_obj_dout_15_rsc_rls_wait_ctrl
    (
  core_wten, dout_15_rsc_rls_obj_iswt0, dout_15_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input dout_15_rsc_rls_obj_iswt0;
  output dout_15_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_15_rsc_rls_obj_ld_core_sct = dout_15_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_dout_15_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_dout_15_rsc_wait_ctrl
    (
  core_wten, dout_15_rsci_iswt0, dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_15_rsci_iswt0;
  output dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_15_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_dout_14_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_dout_14_rsc_wait_ctrl
    (
  core_wten, dout_14_rsci_iswt0, dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_14_rsci_iswt0;
  output dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_14_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_dout_13_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_dout_13_rsc_wait_ctrl
    (
  core_wten, dout_13_rsci_iswt0, dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_13_rsci_iswt0;
  output dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_13_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_dout_12_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_dout_12_rsc_wait_ctrl
    (
  core_wten, dout_12_rsci_iswt0, dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_12_rsci_iswt0;
  output dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_12_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_dout_11_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_dout_11_rsc_wait_ctrl
    (
  core_wten, dout_11_rsci_iswt0, dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_11_rsci_iswt0;
  output dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_11_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_dout_10_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_dout_10_rsc_wait_ctrl
    (
  core_wten, dout_10_rsci_iswt0, dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_10_rsci_iswt0;
  output dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_10_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_dout_9_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_dout_9_rsc_wait_ctrl
    (
  core_wten, dout_9_rsci_iswt0, dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_9_rsci_iswt0;
  output dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_9_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_dout_8_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_dout_8_rsc_wait_ctrl
    (
  core_wten, dout_8_rsci_iswt0, dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_8_rsci_iswt0;
  output dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_8_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_dout_7_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_dout_7_rsc_wait_ctrl
    (
  core_wten, dout_7_rsci_iswt0, dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_7_rsci_iswt0;
  output dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_7_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_dout_6_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_dout_6_rsc_wait_ctrl
    (
  core_wten, dout_6_rsci_iswt0, dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_6_rsci_iswt0;
  output dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_6_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_dout_5_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_dout_5_rsc_wait_ctrl
    (
  core_wten, dout_5_rsci_iswt0, dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_5_rsci_iswt0;
  output dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_5_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_dout_4_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_dout_4_rsc_wait_ctrl
    (
  core_wten, dout_4_rsci_iswt0, dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_4_rsci_iswt0;
  output dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_4_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_dout_3_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_dout_3_rsc_wait_ctrl
    (
  core_wten, dout_3_rsci_iswt0, dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_3_rsci_iswt0;
  output dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_3_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_dout_2_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_dout_2_rsc_wait_ctrl
    (
  core_wten, dout_2_rsci_iswt0, dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_2_rsci_iswt0;
  output dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_2_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_dout_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_dout_1_rsc_wait_ctrl
    (
  core_wten, dout_1_rsci_iswt0, dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_1_rsci_iswt0;
  output dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_1_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_dout_0_rsc_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_dout_0_rsc_wait_ctrl
    (
  core_wten, dout_0_rsci_iswt0, dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct
);
  input core_wten;
  input dout_0_rsci_iswt0;
  output dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct = dout_0_rsci_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci_din_wait_dp
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci_din_wait_dp (
  clk, rst, din_rsci_oswt, din_rsci_wen_comp, din_rsci_d_mxwt, din_rsci_biwt, din_rsci_bdwt,
      din_rsci_d
);
  input clk;
  input rst;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [1023:0] din_rsci_d_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  input [1023:0] din_rsci_d;


  // Interconnect Declarations
  reg din_rsci_bcwt;
  reg [1023:0] din_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_wen_comp = (~ din_rsci_oswt) | din_rsci_biwt | din_rsci_bcwt;
  assign din_rsci_d_mxwt = MUX_v_1024_2_2(din_rsci_d, din_rsci_d_bfwt, din_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsci_bcwt <= 1'b0;
      din_rsci_d_bfwt <= {512'b0 , 512'b0};
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
      din_rsci_d_bfwt <= din_rsci_d_mxwt;
    end
  end

  function [1023:0] MUX_v_1024_2_2;
    input [1023:0] input_0;
    input [1023:0] input_1;
    input [0:0] sel;
    reg [1023:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_1024_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci_din_wait_ctrl
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci_din_wait_ctrl (
  clk, rst, core_wen, din_rsci_oswt, core_wten, din_rsci_biwt, din_rsci_bdwt, din_rsci_ld_core_sct,
      din_rsci_vd
);
  input clk;
  input rst;
  input core_wen;
  input din_rsci_oswt;
  input core_wten;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  output din_rsci_ld_core_sct;
  input din_rsci_vd;


  // Interconnect Declarations
  wire din_rsci_ogwt;
  wire din_rsci_pdswt0;
  reg din_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_pdswt0 = (~ core_wten) & din_rsci_oswt;
  assign din_rsci_biwt = din_rsci_ogwt & din_rsci_vd;
  assign din_rsci_ogwt = din_rsci_pdswt0 | din_rsci_icwt;
  assign din_rsci_bdwt = din_rsci_oswt & core_wen;
  assign din_rsci_ld_core_sct = din_rsci_oswt & din_rsci_ogwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_rsci_icwt <= 1'b0;
    end
    else begin
      din_rsci_icwt <= ~((~(din_rsci_icwt | din_rsci_pdswt0)) | din_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_160_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_160_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_15_and_nl;
  wire din_15_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_15_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_15_and_nl);
  assign din_15_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_15_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_159_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_159_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_14_and_nl;
  wire din_14_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_14_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_14_and_nl);
  assign din_14_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_14_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_158_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_158_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_13_and_nl;
  wire din_13_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_13_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_13_and_nl);
  assign din_13_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_13_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_157_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_157_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_12_and_nl;
  wire din_12_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_12_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_12_and_nl);
  assign din_12_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_12_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_156_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_156_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_11_and_nl;
  wire din_11_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_11_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_11_and_nl);
  assign din_11_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_11_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_155_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_155_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_10_and_nl;
  wire din_10_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_10_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_10_and_nl);
  assign din_10_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_10_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_154_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_154_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_9_and_nl;
  wire din_9_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_9_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_9_and_nl);
  assign din_9_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_9_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_153_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_153_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_8_and_nl;
  wire din_8_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_8_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_8_and_nl);
  assign din_8_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_8_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_152_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_152_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_7_and_nl;
  wire din_7_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_7_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_7_and_nl);
  assign din_7_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_7_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_151_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_151_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_6_and_nl;
  wire din_6_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_6_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_6_and_nl);
  assign din_6_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_6_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_150_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_150_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_5_and_nl;
  wire din_5_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_5_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_5_and_nl);
  assign din_5_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_5_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_149_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_149_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_4_and_nl;
  wire din_4_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_4_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_4_and_nl);
  assign din_4_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_4_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_148_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_148_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_3_and_nl;
  wire din_3_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_3_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_3_and_nl);
  assign din_3_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_3_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_147_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_147_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_2_and_nl;
  wire din_2_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_2_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_2_and_nl);
  assign din_2_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_2_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_146_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_146_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_1_and_nl;
  wire din_1_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_1_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_1_and_nl);
  assign din_1_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_1_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_145_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
// ------------------------------------------------------------------


module catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_145_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
    (
  douta, dinb, addrb, addra, csb_n, csa_n, addra_d, addrb_d, dinb_d, douta_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] douta;
  output [63:0] dinb;
  output [7:0] addrb;
  output [7:0] addra;
  output csb_n;
  output csa_n;
  input [7:0] addra_d;
  input [7:0] addrb_d;
  input [63:0] dinb_d;
  output [63:0] douta_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_0_and_nl;
  wire din_0_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign douta_d = douta;
  assign dinb = (dinb_d);
  assign addrb = (addrb_d);
  assign addra = (addra_d);
  assign din_0_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csa_n = (din_0_and_nl);
  assign din_0_and_1_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb_n = (din_0_and_1_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_staller
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_staller (
  clk, rst, core_wen, core_wten, dout_rsci_wen_comp, din_15_rsc_req_obj_wen_comp,
      din_14_rsc_req_obj_wen_comp, din_13_rsc_req_obj_wen_comp, din_12_rsc_req_obj_wen_comp,
      din_11_rsc_req_obj_wen_comp, din_10_rsc_req_obj_wen_comp, din_9_rsc_req_obj_wen_comp,
      din_8_rsc_req_obj_wen_comp, din_7_rsc_req_obj_wen_comp, din_6_rsc_req_obj_wen_comp,
      din_5_rsc_req_obj_wen_comp, din_4_rsc_req_obj_wen_comp, din_3_rsc_req_obj_wen_comp,
      din_2_rsc_req_obj_wen_comp, din_1_rsc_req_obj_wen_comp, din_0_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input dout_rsci_wen_comp;
  input din_15_rsc_req_obj_wen_comp;
  input din_14_rsc_req_obj_wen_comp;
  input din_13_rsc_req_obj_wen_comp;
  input din_12_rsc_req_obj_wen_comp;
  input din_11_rsc_req_obj_wen_comp;
  input din_10_rsc_req_obj_wen_comp;
  input din_9_rsc_req_obj_wen_comp;
  input din_8_rsc_req_obj_wen_comp;
  input din_7_rsc_req_obj_wen_comp;
  input din_6_rsc_req_obj_wen_comp;
  input din_5_rsc_req_obj_wen_comp;
  input din_4_rsc_req_obj_wen_comp;
  input din_3_rsc_req_obj_wen_comp;
  input din_2_rsc_req_obj_wen_comp;
  input din_1_rsc_req_obj_wen_comp;
  input din_0_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = dout_rsci_wen_comp & din_15_rsc_req_obj_wen_comp & din_14_rsc_req_obj_wen_comp
      & din_13_rsc_req_obj_wen_comp & din_12_rsc_req_obj_wen_comp & din_11_rsc_req_obj_wen_comp
      & din_10_rsc_req_obj_wen_comp & din_9_rsc_req_obj_wen_comp & din_8_rsc_req_obj_wen_comp
      & din_7_rsc_req_obj_wen_comp & din_6_rsc_req_obj_wen_comp & din_5_rsc_req_obj_wen_comp
      & din_4_rsc_req_obj_wen_comp & din_3_rsc_req_obj_wen_comp & din_2_rsc_req_obj_wen_comp
      & din_1_rsc_req_obj_wen_comp & din_0_rsc_req_obj_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj_din_0_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj_din_0_rsc_req_wait_dp
    (
  clk, rst, din_0_rsc_req_obj_oswt, din_0_rsc_req_obj_wen_comp, din_0_rsc_req_obj_biwt,
      din_0_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_0_rsc_req_obj_oswt;
  output din_0_rsc_req_obj_wen_comp;
  input din_0_rsc_req_obj_biwt;
  input din_0_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_0_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_0_rsc_req_obj_wen_comp = (~ din_0_rsc_req_obj_oswt) | din_0_rsc_req_obj_biwt
      | din_0_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_0_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_0_rsc_req_obj_bcwt <= ~((~(din_0_rsc_req_obj_bcwt | din_0_rsc_req_obj_biwt))
          | din_0_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj_din_0_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj_din_0_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_0_rsc_req_obj_oswt, din_0_rsc_req_obj_vd, din_0_rsc_req_obj_biwt,
      din_0_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_0_rsc_req_obj_oswt;
  input din_0_rsc_req_obj_vd;
  output din_0_rsc_req_obj_biwt;
  output din_0_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_0_rsc_req_obj_pdswt0;
  reg din_0_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_0_rsc_req_obj_pdswt0 = (~ core_wten) & din_0_rsc_req_obj_oswt;
  assign din_0_rsc_req_obj_biwt = (din_0_rsc_req_obj_pdswt0 | din_0_rsc_req_obj_icwt)
      & din_0_rsc_req_obj_vd;
  assign din_0_rsc_req_obj_bdwt = din_0_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_0_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_0_rsc_req_obj_icwt <= ~((~(din_0_rsc_req_obj_icwt | din_0_rsc_req_obj_pdswt0))
          | din_0_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj_din_1_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj_din_1_rsc_req_wait_dp
    (
  clk, rst, din_1_rsc_req_obj_oswt, din_1_rsc_req_obj_wen_comp, din_1_rsc_req_obj_biwt,
      din_1_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_1_rsc_req_obj_oswt;
  output din_1_rsc_req_obj_wen_comp;
  input din_1_rsc_req_obj_biwt;
  input din_1_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_1_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_1_rsc_req_obj_wen_comp = (~ din_1_rsc_req_obj_oswt) | din_1_rsc_req_obj_biwt
      | din_1_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_1_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_1_rsc_req_obj_bcwt <= ~((~(din_1_rsc_req_obj_bcwt | din_1_rsc_req_obj_biwt))
          | din_1_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj_din_1_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj_din_1_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_1_rsc_req_obj_oswt, din_1_rsc_req_obj_vd, din_1_rsc_req_obj_biwt,
      din_1_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_1_rsc_req_obj_oswt;
  input din_1_rsc_req_obj_vd;
  output din_1_rsc_req_obj_biwt;
  output din_1_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_1_rsc_req_obj_pdswt0;
  reg din_1_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_1_rsc_req_obj_pdswt0 = (~ core_wten) & din_1_rsc_req_obj_oswt;
  assign din_1_rsc_req_obj_biwt = (din_1_rsc_req_obj_pdswt0 | din_1_rsc_req_obj_icwt)
      & din_1_rsc_req_obj_vd;
  assign din_1_rsc_req_obj_bdwt = din_1_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_1_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_1_rsc_req_obj_icwt <= ~((~(din_1_rsc_req_obj_icwt | din_1_rsc_req_obj_pdswt0))
          | din_1_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj_din_2_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj_din_2_rsc_req_wait_dp
    (
  clk, rst, din_2_rsc_req_obj_oswt, din_2_rsc_req_obj_wen_comp, din_2_rsc_req_obj_biwt,
      din_2_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_2_rsc_req_obj_oswt;
  output din_2_rsc_req_obj_wen_comp;
  input din_2_rsc_req_obj_biwt;
  input din_2_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_2_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_2_rsc_req_obj_wen_comp = (~ din_2_rsc_req_obj_oswt) | din_2_rsc_req_obj_biwt
      | din_2_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_2_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_2_rsc_req_obj_bcwt <= ~((~(din_2_rsc_req_obj_bcwt | din_2_rsc_req_obj_biwt))
          | din_2_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj_din_2_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj_din_2_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_2_rsc_req_obj_oswt, din_2_rsc_req_obj_vd, din_2_rsc_req_obj_biwt,
      din_2_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_2_rsc_req_obj_oswt;
  input din_2_rsc_req_obj_vd;
  output din_2_rsc_req_obj_biwt;
  output din_2_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_2_rsc_req_obj_pdswt0;
  reg din_2_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_2_rsc_req_obj_pdswt0 = (~ core_wten) & din_2_rsc_req_obj_oswt;
  assign din_2_rsc_req_obj_biwt = (din_2_rsc_req_obj_pdswt0 | din_2_rsc_req_obj_icwt)
      & din_2_rsc_req_obj_vd;
  assign din_2_rsc_req_obj_bdwt = din_2_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_2_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_2_rsc_req_obj_icwt <= ~((~(din_2_rsc_req_obj_icwt | din_2_rsc_req_obj_pdswt0))
          | din_2_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj_din_3_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj_din_3_rsc_req_wait_dp
    (
  clk, rst, din_3_rsc_req_obj_oswt, din_3_rsc_req_obj_wen_comp, din_3_rsc_req_obj_biwt,
      din_3_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_3_rsc_req_obj_oswt;
  output din_3_rsc_req_obj_wen_comp;
  input din_3_rsc_req_obj_biwt;
  input din_3_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_3_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_3_rsc_req_obj_wen_comp = (~ din_3_rsc_req_obj_oswt) | din_3_rsc_req_obj_biwt
      | din_3_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_3_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_3_rsc_req_obj_bcwt <= ~((~(din_3_rsc_req_obj_bcwt | din_3_rsc_req_obj_biwt))
          | din_3_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj_din_3_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj_din_3_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_3_rsc_req_obj_oswt, din_3_rsc_req_obj_vd, din_3_rsc_req_obj_biwt,
      din_3_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_3_rsc_req_obj_oswt;
  input din_3_rsc_req_obj_vd;
  output din_3_rsc_req_obj_biwt;
  output din_3_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_3_rsc_req_obj_pdswt0;
  reg din_3_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_3_rsc_req_obj_pdswt0 = (~ core_wten) & din_3_rsc_req_obj_oswt;
  assign din_3_rsc_req_obj_biwt = (din_3_rsc_req_obj_pdswt0 | din_3_rsc_req_obj_icwt)
      & din_3_rsc_req_obj_vd;
  assign din_3_rsc_req_obj_bdwt = din_3_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_3_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_3_rsc_req_obj_icwt <= ~((~(din_3_rsc_req_obj_icwt | din_3_rsc_req_obj_pdswt0))
          | din_3_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj_din_4_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj_din_4_rsc_req_wait_dp
    (
  clk, rst, din_4_rsc_req_obj_oswt, din_4_rsc_req_obj_wen_comp, din_4_rsc_req_obj_biwt,
      din_4_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_4_rsc_req_obj_oswt;
  output din_4_rsc_req_obj_wen_comp;
  input din_4_rsc_req_obj_biwt;
  input din_4_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_4_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_4_rsc_req_obj_wen_comp = (~ din_4_rsc_req_obj_oswt) | din_4_rsc_req_obj_biwt
      | din_4_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_4_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_4_rsc_req_obj_bcwt <= ~((~(din_4_rsc_req_obj_bcwt | din_4_rsc_req_obj_biwt))
          | din_4_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj_din_4_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj_din_4_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_4_rsc_req_obj_oswt, din_4_rsc_req_obj_vd, din_4_rsc_req_obj_biwt,
      din_4_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_4_rsc_req_obj_oswt;
  input din_4_rsc_req_obj_vd;
  output din_4_rsc_req_obj_biwt;
  output din_4_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_4_rsc_req_obj_pdswt0;
  reg din_4_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_4_rsc_req_obj_pdswt0 = (~ core_wten) & din_4_rsc_req_obj_oswt;
  assign din_4_rsc_req_obj_biwt = (din_4_rsc_req_obj_pdswt0 | din_4_rsc_req_obj_icwt)
      & din_4_rsc_req_obj_vd;
  assign din_4_rsc_req_obj_bdwt = din_4_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_4_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_4_rsc_req_obj_icwt <= ~((~(din_4_rsc_req_obj_icwt | din_4_rsc_req_obj_pdswt0))
          | din_4_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj_din_5_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj_din_5_rsc_req_wait_dp
    (
  clk, rst, din_5_rsc_req_obj_oswt, din_5_rsc_req_obj_wen_comp, din_5_rsc_req_obj_biwt,
      din_5_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_5_rsc_req_obj_oswt;
  output din_5_rsc_req_obj_wen_comp;
  input din_5_rsc_req_obj_biwt;
  input din_5_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_5_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_5_rsc_req_obj_wen_comp = (~ din_5_rsc_req_obj_oswt) | din_5_rsc_req_obj_biwt
      | din_5_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_5_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_5_rsc_req_obj_bcwt <= ~((~(din_5_rsc_req_obj_bcwt | din_5_rsc_req_obj_biwt))
          | din_5_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj_din_5_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj_din_5_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_5_rsc_req_obj_oswt, din_5_rsc_req_obj_vd, din_5_rsc_req_obj_biwt,
      din_5_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_5_rsc_req_obj_oswt;
  input din_5_rsc_req_obj_vd;
  output din_5_rsc_req_obj_biwt;
  output din_5_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_5_rsc_req_obj_pdswt0;
  reg din_5_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_5_rsc_req_obj_pdswt0 = (~ core_wten) & din_5_rsc_req_obj_oswt;
  assign din_5_rsc_req_obj_biwt = (din_5_rsc_req_obj_pdswt0 | din_5_rsc_req_obj_icwt)
      & din_5_rsc_req_obj_vd;
  assign din_5_rsc_req_obj_bdwt = din_5_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_5_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_5_rsc_req_obj_icwt <= ~((~(din_5_rsc_req_obj_icwt | din_5_rsc_req_obj_pdswt0))
          | din_5_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj_din_6_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj_din_6_rsc_req_wait_dp
    (
  clk, rst, din_6_rsc_req_obj_oswt, din_6_rsc_req_obj_wen_comp, din_6_rsc_req_obj_biwt,
      din_6_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_6_rsc_req_obj_oswt;
  output din_6_rsc_req_obj_wen_comp;
  input din_6_rsc_req_obj_biwt;
  input din_6_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_6_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_6_rsc_req_obj_wen_comp = (~ din_6_rsc_req_obj_oswt) | din_6_rsc_req_obj_biwt
      | din_6_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_6_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_6_rsc_req_obj_bcwt <= ~((~(din_6_rsc_req_obj_bcwt | din_6_rsc_req_obj_biwt))
          | din_6_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj_din_6_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj_din_6_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_6_rsc_req_obj_oswt, din_6_rsc_req_obj_vd, din_6_rsc_req_obj_biwt,
      din_6_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_6_rsc_req_obj_oswt;
  input din_6_rsc_req_obj_vd;
  output din_6_rsc_req_obj_biwt;
  output din_6_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_6_rsc_req_obj_pdswt0;
  reg din_6_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_6_rsc_req_obj_pdswt0 = (~ core_wten) & din_6_rsc_req_obj_oswt;
  assign din_6_rsc_req_obj_biwt = (din_6_rsc_req_obj_pdswt0 | din_6_rsc_req_obj_icwt)
      & din_6_rsc_req_obj_vd;
  assign din_6_rsc_req_obj_bdwt = din_6_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_6_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_6_rsc_req_obj_icwt <= ~((~(din_6_rsc_req_obj_icwt | din_6_rsc_req_obj_pdswt0))
          | din_6_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj_din_7_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj_din_7_rsc_req_wait_dp
    (
  clk, rst, din_7_rsc_req_obj_oswt, din_7_rsc_req_obj_wen_comp, din_7_rsc_req_obj_biwt,
      din_7_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_7_rsc_req_obj_oswt;
  output din_7_rsc_req_obj_wen_comp;
  input din_7_rsc_req_obj_biwt;
  input din_7_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_7_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_7_rsc_req_obj_wen_comp = (~ din_7_rsc_req_obj_oswt) | din_7_rsc_req_obj_biwt
      | din_7_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_7_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_7_rsc_req_obj_bcwt <= ~((~(din_7_rsc_req_obj_bcwt | din_7_rsc_req_obj_biwt))
          | din_7_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj_din_7_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj_din_7_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_7_rsc_req_obj_oswt, din_7_rsc_req_obj_vd, din_7_rsc_req_obj_biwt,
      din_7_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_7_rsc_req_obj_oswt;
  input din_7_rsc_req_obj_vd;
  output din_7_rsc_req_obj_biwt;
  output din_7_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_7_rsc_req_obj_pdswt0;
  reg din_7_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_7_rsc_req_obj_pdswt0 = (~ core_wten) & din_7_rsc_req_obj_oswt;
  assign din_7_rsc_req_obj_biwt = (din_7_rsc_req_obj_pdswt0 | din_7_rsc_req_obj_icwt)
      & din_7_rsc_req_obj_vd;
  assign din_7_rsc_req_obj_bdwt = din_7_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_7_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_7_rsc_req_obj_icwt <= ~((~(din_7_rsc_req_obj_icwt | din_7_rsc_req_obj_pdswt0))
          | din_7_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj_din_8_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj_din_8_rsc_req_wait_dp
    (
  clk, rst, din_8_rsc_req_obj_oswt, din_8_rsc_req_obj_wen_comp, din_8_rsc_req_obj_biwt,
      din_8_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_8_rsc_req_obj_oswt;
  output din_8_rsc_req_obj_wen_comp;
  input din_8_rsc_req_obj_biwt;
  input din_8_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_8_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_8_rsc_req_obj_wen_comp = (~ din_8_rsc_req_obj_oswt) | din_8_rsc_req_obj_biwt
      | din_8_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_8_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_8_rsc_req_obj_bcwt <= ~((~(din_8_rsc_req_obj_bcwt | din_8_rsc_req_obj_biwt))
          | din_8_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj_din_8_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj_din_8_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_8_rsc_req_obj_oswt, din_8_rsc_req_obj_vd, din_8_rsc_req_obj_biwt,
      din_8_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_8_rsc_req_obj_oswt;
  input din_8_rsc_req_obj_vd;
  output din_8_rsc_req_obj_biwt;
  output din_8_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_8_rsc_req_obj_pdswt0;
  reg din_8_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_8_rsc_req_obj_pdswt0 = (~ core_wten) & din_8_rsc_req_obj_oswt;
  assign din_8_rsc_req_obj_biwt = (din_8_rsc_req_obj_pdswt0 | din_8_rsc_req_obj_icwt)
      & din_8_rsc_req_obj_vd;
  assign din_8_rsc_req_obj_bdwt = din_8_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_8_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_8_rsc_req_obj_icwt <= ~((~(din_8_rsc_req_obj_icwt | din_8_rsc_req_obj_pdswt0))
          | din_8_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj_din_9_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj_din_9_rsc_req_wait_dp
    (
  clk, rst, din_9_rsc_req_obj_oswt, din_9_rsc_req_obj_wen_comp, din_9_rsc_req_obj_biwt,
      din_9_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_9_rsc_req_obj_oswt;
  output din_9_rsc_req_obj_wen_comp;
  input din_9_rsc_req_obj_biwt;
  input din_9_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_9_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_9_rsc_req_obj_wen_comp = (~ din_9_rsc_req_obj_oswt) | din_9_rsc_req_obj_biwt
      | din_9_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_9_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_9_rsc_req_obj_bcwt <= ~((~(din_9_rsc_req_obj_bcwt | din_9_rsc_req_obj_biwt))
          | din_9_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj_din_9_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj_din_9_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_9_rsc_req_obj_oswt, din_9_rsc_req_obj_vd, din_9_rsc_req_obj_biwt,
      din_9_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_9_rsc_req_obj_oswt;
  input din_9_rsc_req_obj_vd;
  output din_9_rsc_req_obj_biwt;
  output din_9_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_9_rsc_req_obj_pdswt0;
  reg din_9_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_9_rsc_req_obj_pdswt0 = (~ core_wten) & din_9_rsc_req_obj_oswt;
  assign din_9_rsc_req_obj_biwt = (din_9_rsc_req_obj_pdswt0 | din_9_rsc_req_obj_icwt)
      & din_9_rsc_req_obj_vd;
  assign din_9_rsc_req_obj_bdwt = din_9_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_9_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_9_rsc_req_obj_icwt <= ~((~(din_9_rsc_req_obj_icwt | din_9_rsc_req_obj_pdswt0))
          | din_9_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj_din_10_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj_din_10_rsc_req_wait_dp
    (
  clk, rst, din_10_rsc_req_obj_oswt, din_10_rsc_req_obj_wen_comp, din_10_rsc_req_obj_biwt,
      din_10_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_10_rsc_req_obj_oswt;
  output din_10_rsc_req_obj_wen_comp;
  input din_10_rsc_req_obj_biwt;
  input din_10_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_10_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_10_rsc_req_obj_wen_comp = (~ din_10_rsc_req_obj_oswt) | din_10_rsc_req_obj_biwt
      | din_10_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_10_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_10_rsc_req_obj_bcwt <= ~((~(din_10_rsc_req_obj_bcwt | din_10_rsc_req_obj_biwt))
          | din_10_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj_din_10_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj_din_10_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_10_rsc_req_obj_oswt, din_10_rsc_req_obj_vd,
      din_10_rsc_req_obj_biwt, din_10_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_10_rsc_req_obj_oswt;
  input din_10_rsc_req_obj_vd;
  output din_10_rsc_req_obj_biwt;
  output din_10_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_10_rsc_req_obj_pdswt0;
  reg din_10_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_10_rsc_req_obj_pdswt0 = (~ core_wten) & din_10_rsc_req_obj_oswt;
  assign din_10_rsc_req_obj_biwt = (din_10_rsc_req_obj_pdswt0 | din_10_rsc_req_obj_icwt)
      & din_10_rsc_req_obj_vd;
  assign din_10_rsc_req_obj_bdwt = din_10_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_10_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_10_rsc_req_obj_icwt <= ~((~(din_10_rsc_req_obj_icwt | din_10_rsc_req_obj_pdswt0))
          | din_10_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj_din_11_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj_din_11_rsc_req_wait_dp
    (
  clk, rst, din_11_rsc_req_obj_oswt, din_11_rsc_req_obj_wen_comp, din_11_rsc_req_obj_biwt,
      din_11_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_11_rsc_req_obj_oswt;
  output din_11_rsc_req_obj_wen_comp;
  input din_11_rsc_req_obj_biwt;
  input din_11_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_11_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_11_rsc_req_obj_wen_comp = (~ din_11_rsc_req_obj_oswt) | din_11_rsc_req_obj_biwt
      | din_11_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_11_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_11_rsc_req_obj_bcwt <= ~((~(din_11_rsc_req_obj_bcwt | din_11_rsc_req_obj_biwt))
          | din_11_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj_din_11_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj_din_11_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_11_rsc_req_obj_oswt, din_11_rsc_req_obj_vd,
      din_11_rsc_req_obj_biwt, din_11_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_11_rsc_req_obj_oswt;
  input din_11_rsc_req_obj_vd;
  output din_11_rsc_req_obj_biwt;
  output din_11_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_11_rsc_req_obj_pdswt0;
  reg din_11_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_11_rsc_req_obj_pdswt0 = (~ core_wten) & din_11_rsc_req_obj_oswt;
  assign din_11_rsc_req_obj_biwt = (din_11_rsc_req_obj_pdswt0 | din_11_rsc_req_obj_icwt)
      & din_11_rsc_req_obj_vd;
  assign din_11_rsc_req_obj_bdwt = din_11_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_11_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_11_rsc_req_obj_icwt <= ~((~(din_11_rsc_req_obj_icwt | din_11_rsc_req_obj_pdswt0))
          | din_11_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj_din_12_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj_din_12_rsc_req_wait_dp
    (
  clk, rst, din_12_rsc_req_obj_oswt, din_12_rsc_req_obj_wen_comp, din_12_rsc_req_obj_biwt,
      din_12_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_12_rsc_req_obj_oswt;
  output din_12_rsc_req_obj_wen_comp;
  input din_12_rsc_req_obj_biwt;
  input din_12_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_12_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_12_rsc_req_obj_wen_comp = (~ din_12_rsc_req_obj_oswt) | din_12_rsc_req_obj_biwt
      | din_12_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_12_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_12_rsc_req_obj_bcwt <= ~((~(din_12_rsc_req_obj_bcwt | din_12_rsc_req_obj_biwt))
          | din_12_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj_din_12_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj_din_12_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_12_rsc_req_obj_oswt, din_12_rsc_req_obj_vd,
      din_12_rsc_req_obj_biwt, din_12_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_12_rsc_req_obj_oswt;
  input din_12_rsc_req_obj_vd;
  output din_12_rsc_req_obj_biwt;
  output din_12_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_12_rsc_req_obj_pdswt0;
  reg din_12_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_12_rsc_req_obj_pdswt0 = (~ core_wten) & din_12_rsc_req_obj_oswt;
  assign din_12_rsc_req_obj_biwt = (din_12_rsc_req_obj_pdswt0 | din_12_rsc_req_obj_icwt)
      & din_12_rsc_req_obj_vd;
  assign din_12_rsc_req_obj_bdwt = din_12_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_12_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_12_rsc_req_obj_icwt <= ~((~(din_12_rsc_req_obj_icwt | din_12_rsc_req_obj_pdswt0))
          | din_12_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj_din_13_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj_din_13_rsc_req_wait_dp
    (
  clk, rst, din_13_rsc_req_obj_oswt, din_13_rsc_req_obj_wen_comp, din_13_rsc_req_obj_biwt,
      din_13_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_13_rsc_req_obj_oswt;
  output din_13_rsc_req_obj_wen_comp;
  input din_13_rsc_req_obj_biwt;
  input din_13_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_13_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_13_rsc_req_obj_wen_comp = (~ din_13_rsc_req_obj_oswt) | din_13_rsc_req_obj_biwt
      | din_13_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_13_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_13_rsc_req_obj_bcwt <= ~((~(din_13_rsc_req_obj_bcwt | din_13_rsc_req_obj_biwt))
          | din_13_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj_din_13_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj_din_13_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_13_rsc_req_obj_oswt, din_13_rsc_req_obj_vd,
      din_13_rsc_req_obj_biwt, din_13_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_13_rsc_req_obj_oswt;
  input din_13_rsc_req_obj_vd;
  output din_13_rsc_req_obj_biwt;
  output din_13_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_13_rsc_req_obj_pdswt0;
  reg din_13_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_13_rsc_req_obj_pdswt0 = (~ core_wten) & din_13_rsc_req_obj_oswt;
  assign din_13_rsc_req_obj_biwt = (din_13_rsc_req_obj_pdswt0 | din_13_rsc_req_obj_icwt)
      & din_13_rsc_req_obj_vd;
  assign din_13_rsc_req_obj_bdwt = din_13_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_13_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_13_rsc_req_obj_icwt <= ~((~(din_13_rsc_req_obj_icwt | din_13_rsc_req_obj_pdswt0))
          | din_13_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj_din_14_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj_din_14_rsc_req_wait_dp
    (
  clk, rst, din_14_rsc_req_obj_oswt, din_14_rsc_req_obj_wen_comp, din_14_rsc_req_obj_biwt,
      din_14_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_14_rsc_req_obj_oswt;
  output din_14_rsc_req_obj_wen_comp;
  input din_14_rsc_req_obj_biwt;
  input din_14_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_14_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_14_rsc_req_obj_wen_comp = (~ din_14_rsc_req_obj_oswt) | din_14_rsc_req_obj_biwt
      | din_14_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_14_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_14_rsc_req_obj_bcwt <= ~((~(din_14_rsc_req_obj_bcwt | din_14_rsc_req_obj_biwt))
          | din_14_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj_din_14_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj_din_14_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_14_rsc_req_obj_oswt, din_14_rsc_req_obj_vd,
      din_14_rsc_req_obj_biwt, din_14_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_14_rsc_req_obj_oswt;
  input din_14_rsc_req_obj_vd;
  output din_14_rsc_req_obj_biwt;
  output din_14_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_14_rsc_req_obj_pdswt0;
  reg din_14_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_14_rsc_req_obj_pdswt0 = (~ core_wten) & din_14_rsc_req_obj_oswt;
  assign din_14_rsc_req_obj_biwt = (din_14_rsc_req_obj_pdswt0 | din_14_rsc_req_obj_icwt)
      & din_14_rsc_req_obj_vd;
  assign din_14_rsc_req_obj_bdwt = din_14_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_14_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_14_rsc_req_obj_icwt <= ~((~(din_14_rsc_req_obj_icwt | din_14_rsc_req_obj_pdswt0))
          | din_14_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj_din_15_rsc_req_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj_din_15_rsc_req_wait_dp
    (
  clk, rst, din_15_rsc_req_obj_oswt, din_15_rsc_req_obj_wen_comp, din_15_rsc_req_obj_biwt,
      din_15_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input din_15_rsc_req_obj_oswt;
  output din_15_rsc_req_obj_wen_comp;
  input din_15_rsc_req_obj_biwt;
  input din_15_rsc_req_obj_bdwt;


  // Interconnect Declarations
  reg din_15_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_15_rsc_req_obj_wen_comp = (~ din_15_rsc_req_obj_oswt) | din_15_rsc_req_obj_biwt
      | din_15_rsc_req_obj_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      din_15_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_15_rsc_req_obj_bcwt <= ~((~(din_15_rsc_req_obj_bcwt | din_15_rsc_req_obj_biwt))
          | din_15_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj_din_15_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj_din_15_rsc_req_wait_ctrl
    (
  clk, rst, core_wen, core_wten, din_15_rsc_req_obj_oswt, din_15_rsc_req_obj_vd,
      din_15_rsc_req_obj_biwt, din_15_rsc_req_obj_bdwt
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input din_15_rsc_req_obj_oswt;
  input din_15_rsc_req_obj_vd;
  output din_15_rsc_req_obj_biwt;
  output din_15_rsc_req_obj_bdwt;


  // Interconnect Declarations
  wire din_15_rsc_req_obj_pdswt0;
  reg din_15_rsc_req_obj_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_15_rsc_req_obj_pdswt0 = (~ core_wten) & din_15_rsc_req_obj_oswt;
  assign din_15_rsc_req_obj_biwt = (din_15_rsc_req_obj_pdswt0 | din_15_rsc_req_obj_icwt)
      & din_15_rsc_req_obj_vd;
  assign din_15_rsc_req_obj_bdwt = din_15_rsc_req_obj_oswt & core_wen;
  always @(posedge clk) begin
    if ( rst ) begin
      din_15_rsc_req_obj_icwt <= 1'b0;
    end
    else begin
      din_15_rsc_req_obj_icwt <= ~((~(din_15_rsc_req_obj_icwt | din_15_rsc_req_obj_pdswt0))
          | din_15_rsc_req_obj_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_rls_obj_din_15_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_rls_obj_din_15_rsc_rls_wait_ctrl
    (
  core_wten, din_15_rsc_rls_obj_iswt0, din_15_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_15_rsc_rls_obj_iswt0;
  output din_15_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_15_rsc_rls_obj_ld_core_sct = din_15_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_rls_obj_din_14_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_rls_obj_din_14_rsc_rls_wait_ctrl
    (
  core_wten, din_14_rsc_rls_obj_iswt0, din_14_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_14_rsc_rls_obj_iswt0;
  output din_14_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_14_rsc_rls_obj_ld_core_sct = din_14_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_rls_obj_din_13_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_rls_obj_din_13_rsc_rls_wait_ctrl
    (
  core_wten, din_13_rsc_rls_obj_iswt0, din_13_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_13_rsc_rls_obj_iswt0;
  output din_13_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_13_rsc_rls_obj_ld_core_sct = din_13_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_rls_obj_din_12_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_rls_obj_din_12_rsc_rls_wait_ctrl
    (
  core_wten, din_12_rsc_rls_obj_iswt0, din_12_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_12_rsc_rls_obj_iswt0;
  output din_12_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_12_rsc_rls_obj_ld_core_sct = din_12_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_rls_obj_din_11_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_rls_obj_din_11_rsc_rls_wait_ctrl
    (
  core_wten, din_11_rsc_rls_obj_iswt0, din_11_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_11_rsc_rls_obj_iswt0;
  output din_11_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_11_rsc_rls_obj_ld_core_sct = din_11_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_rls_obj_din_10_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_rls_obj_din_10_rsc_rls_wait_ctrl
    (
  core_wten, din_10_rsc_rls_obj_iswt0, din_10_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_10_rsc_rls_obj_iswt0;
  output din_10_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_10_rsc_rls_obj_ld_core_sct = din_10_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_rls_obj_din_9_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_rls_obj_din_9_rsc_rls_wait_ctrl
    (
  core_wten, din_9_rsc_rls_obj_iswt0, din_9_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_9_rsc_rls_obj_iswt0;
  output din_9_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_9_rsc_rls_obj_ld_core_sct = din_9_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_rls_obj_din_8_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_rls_obj_din_8_rsc_rls_wait_ctrl
    (
  core_wten, din_8_rsc_rls_obj_iswt0, din_8_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_8_rsc_rls_obj_iswt0;
  output din_8_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_8_rsc_rls_obj_ld_core_sct = din_8_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_rls_obj_din_7_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_rls_obj_din_7_rsc_rls_wait_ctrl
    (
  core_wten, din_7_rsc_rls_obj_iswt0, din_7_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_7_rsc_rls_obj_iswt0;
  output din_7_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_7_rsc_rls_obj_ld_core_sct = din_7_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_rls_obj_din_6_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_rls_obj_din_6_rsc_rls_wait_ctrl
    (
  core_wten, din_6_rsc_rls_obj_iswt0, din_6_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_6_rsc_rls_obj_iswt0;
  output din_6_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_6_rsc_rls_obj_ld_core_sct = din_6_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_rls_obj_din_5_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_rls_obj_din_5_rsc_rls_wait_ctrl
    (
  core_wten, din_5_rsc_rls_obj_iswt0, din_5_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_5_rsc_rls_obj_iswt0;
  output din_5_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_5_rsc_rls_obj_ld_core_sct = din_5_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_rls_obj_din_4_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_rls_obj_din_4_rsc_rls_wait_ctrl
    (
  core_wten, din_4_rsc_rls_obj_iswt0, din_4_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_4_rsc_rls_obj_iswt0;
  output din_4_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_4_rsc_rls_obj_ld_core_sct = din_4_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_rls_obj_din_3_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_rls_obj_din_3_rsc_rls_wait_ctrl
    (
  core_wten, din_3_rsc_rls_obj_iswt0, din_3_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_3_rsc_rls_obj_iswt0;
  output din_3_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_3_rsc_rls_obj_ld_core_sct = din_3_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_rls_obj_din_2_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_rls_obj_din_2_rsc_rls_wait_ctrl
    (
  core_wten, din_2_rsc_rls_obj_iswt0, din_2_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_2_rsc_rls_obj_iswt0;
  output din_2_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_2_rsc_rls_obj_ld_core_sct = din_2_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_rls_obj_din_1_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_rls_obj_din_1_rsc_rls_wait_ctrl
    (
  core_wten, din_1_rsc_rls_obj_iswt0, din_1_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_1_rsc_rls_obj_iswt0;
  output din_1_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_1_rsc_rls_obj_ld_core_sct = din_1_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_rls_obj_din_0_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_rls_obj_din_0_rsc_rls_wait_ctrl
    (
  core_wten, din_0_rsc_rls_obj_iswt0, din_0_rsc_rls_obj_ld_core_sct
);
  input core_wten;
  input din_0_rsc_rls_obj_iswt0;
  output din_0_rsc_rls_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_0_rsc_rls_obj_ld_core_sct = din_0_rsc_rls_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_dout_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_dout_wait_dp (
  clk, rst, dout_rsci_oswt, dout_rsci_wen_comp, dout_rsci_biwt, dout_rsci_bdwt
);
  input clk;
  input rst;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input dout_rsci_biwt;
  input dout_rsci_bdwt;


  // Interconnect Declarations
  reg dout_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_wen_comp = (~ dout_rsci_oswt) | dout_rsci_biwt | dout_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_bcwt <= 1'b0;
    end
    else begin
      dout_rsci_bcwt <= ~((~(dout_rsci_bcwt | dout_rsci_biwt)) | dout_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_dout_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_dout_wait_ctrl (
  clk, rst, core_wen, core_wten, dout_rsci_oswt, dout_rsci_biwt, dout_rsci_bdwt,
      dout_rsci_ld_core_sct, dout_rsci_vd
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input dout_rsci_oswt;
  output dout_rsci_biwt;
  output dout_rsci_bdwt;
  output dout_rsci_ld_core_sct;
  input dout_rsci_vd;


  // Interconnect Declarations
  wire dout_rsci_ogwt;
  wire dout_rsci_pdswt0;
  reg dout_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_pdswt0 = (~ core_wten) & dout_rsci_oswt;
  assign dout_rsci_biwt = dout_rsci_ogwt & dout_rsci_vd;
  assign dout_rsci_ogwt = dout_rsci_pdswt0 | dout_rsci_icwt;
  assign dout_rsci_bdwt = dout_rsci_oswt & core_wen;
  assign dout_rsci_ld_core_sct = dout_rsci_oswt & dout_rsci_ogwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_icwt <= 1'b0;
    end
    else begin
      dout_rsci_icwt <= ~((~(dout_rsci_icwt | dout_rsci_pdswt0)) | dout_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_din_15_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_din_15_rsc_wait_dp (
  clk, rst, din_15_rsci_douta_d, din_15_rsci_douta_d_mxwt, din_15_rsci_biwt, din_15_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_15_rsci_douta_d;
  output [63:0] din_15_rsci_douta_d_mxwt;
  input din_15_rsci_biwt;
  input din_15_rsci_bdwt;


  // Interconnect Declarations
  reg din_15_rsci_bcwt;
  reg [63:0] din_15_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_15_rsci_douta_d_mxwt = MUX_v_64_2_2(din_15_rsci_douta_d, din_15_rsci_douta_d_bfwt,
      din_15_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_15_rsci_bcwt <= 1'b0;
      din_15_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_15_rsci_bcwt <= ~((~(din_15_rsci_bcwt | din_15_rsci_biwt)) | din_15_rsci_bdwt);
      din_15_rsci_douta_d_bfwt <= din_15_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_din_15_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_din_15_rsc_wait_ctrl
    (
  core_wen, core_wten, din_15_rsci_oswt, din_15_rsci_biwt, din_15_rsci_bdwt, din_15_rsci_biwt_pff,
      din_15_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_15_rsci_oswt;
  output din_15_rsci_biwt;
  output din_15_rsci_bdwt;
  output din_15_rsci_biwt_pff;
  input din_15_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_15_rsci_bdwt = din_15_rsci_oswt & core_wen;
  assign din_15_rsci_biwt = (~ core_wten) & din_15_rsci_oswt;
  assign din_15_rsci_biwt_pff = core_wen & din_15_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_din_14_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_din_14_rsc_wait_dp (
  clk, rst, din_14_rsci_douta_d, din_14_rsci_douta_d_mxwt, din_14_rsci_biwt, din_14_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_14_rsci_douta_d;
  output [63:0] din_14_rsci_douta_d_mxwt;
  input din_14_rsci_biwt;
  input din_14_rsci_bdwt;


  // Interconnect Declarations
  reg din_14_rsci_bcwt;
  reg [63:0] din_14_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_14_rsci_douta_d_mxwt = MUX_v_64_2_2(din_14_rsci_douta_d, din_14_rsci_douta_d_bfwt,
      din_14_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_14_rsci_bcwt <= 1'b0;
      din_14_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_14_rsci_bcwt <= ~((~(din_14_rsci_bcwt | din_14_rsci_biwt)) | din_14_rsci_bdwt);
      din_14_rsci_douta_d_bfwt <= din_14_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_din_14_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_din_14_rsc_wait_ctrl
    (
  core_wen, core_wten, din_14_rsci_oswt, din_14_rsci_biwt, din_14_rsci_bdwt, din_14_rsci_biwt_pff,
      din_14_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_14_rsci_oswt;
  output din_14_rsci_biwt;
  output din_14_rsci_bdwt;
  output din_14_rsci_biwt_pff;
  input din_14_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_14_rsci_bdwt = din_14_rsci_oswt & core_wen;
  assign din_14_rsci_biwt = (~ core_wten) & din_14_rsci_oswt;
  assign din_14_rsci_biwt_pff = core_wen & din_14_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_din_13_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_din_13_rsc_wait_dp (
  clk, rst, din_13_rsci_douta_d, din_13_rsci_douta_d_mxwt, din_13_rsci_biwt, din_13_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_13_rsci_douta_d;
  output [63:0] din_13_rsci_douta_d_mxwt;
  input din_13_rsci_biwt;
  input din_13_rsci_bdwt;


  // Interconnect Declarations
  reg din_13_rsci_bcwt;
  reg [63:0] din_13_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_13_rsci_douta_d_mxwt = MUX_v_64_2_2(din_13_rsci_douta_d, din_13_rsci_douta_d_bfwt,
      din_13_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_13_rsci_bcwt <= 1'b0;
      din_13_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_13_rsci_bcwt <= ~((~(din_13_rsci_bcwt | din_13_rsci_biwt)) | din_13_rsci_bdwt);
      din_13_rsci_douta_d_bfwt <= din_13_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_din_13_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_din_13_rsc_wait_ctrl
    (
  core_wen, core_wten, din_13_rsci_oswt, din_13_rsci_biwt, din_13_rsci_bdwt, din_13_rsci_biwt_pff,
      din_13_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_13_rsci_oswt;
  output din_13_rsci_biwt;
  output din_13_rsci_bdwt;
  output din_13_rsci_biwt_pff;
  input din_13_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_13_rsci_bdwt = din_13_rsci_oswt & core_wen;
  assign din_13_rsci_biwt = (~ core_wten) & din_13_rsci_oswt;
  assign din_13_rsci_biwt_pff = core_wen & din_13_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_din_12_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_din_12_rsc_wait_dp (
  clk, rst, din_12_rsci_douta_d, din_12_rsci_douta_d_mxwt, din_12_rsci_biwt, din_12_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_12_rsci_douta_d;
  output [63:0] din_12_rsci_douta_d_mxwt;
  input din_12_rsci_biwt;
  input din_12_rsci_bdwt;


  // Interconnect Declarations
  reg din_12_rsci_bcwt;
  reg [63:0] din_12_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_12_rsci_douta_d_mxwt = MUX_v_64_2_2(din_12_rsci_douta_d, din_12_rsci_douta_d_bfwt,
      din_12_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_12_rsci_bcwt <= 1'b0;
      din_12_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_12_rsci_bcwt <= ~((~(din_12_rsci_bcwt | din_12_rsci_biwt)) | din_12_rsci_bdwt);
      din_12_rsci_douta_d_bfwt <= din_12_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_din_12_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_din_12_rsc_wait_ctrl
    (
  core_wen, core_wten, din_12_rsci_oswt, din_12_rsci_biwt, din_12_rsci_bdwt, din_12_rsci_biwt_pff,
      din_12_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_12_rsci_oswt;
  output din_12_rsci_biwt;
  output din_12_rsci_bdwt;
  output din_12_rsci_biwt_pff;
  input din_12_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_12_rsci_bdwt = din_12_rsci_oswt & core_wen;
  assign din_12_rsci_biwt = (~ core_wten) & din_12_rsci_oswt;
  assign din_12_rsci_biwt_pff = core_wen & din_12_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_din_11_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_din_11_rsc_wait_dp (
  clk, rst, din_11_rsci_douta_d, din_11_rsci_douta_d_mxwt, din_11_rsci_biwt, din_11_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_11_rsci_douta_d;
  output [63:0] din_11_rsci_douta_d_mxwt;
  input din_11_rsci_biwt;
  input din_11_rsci_bdwt;


  // Interconnect Declarations
  reg din_11_rsci_bcwt;
  reg [63:0] din_11_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_11_rsci_douta_d_mxwt = MUX_v_64_2_2(din_11_rsci_douta_d, din_11_rsci_douta_d_bfwt,
      din_11_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_11_rsci_bcwt <= 1'b0;
      din_11_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_11_rsci_bcwt <= ~((~(din_11_rsci_bcwt | din_11_rsci_biwt)) | din_11_rsci_bdwt);
      din_11_rsci_douta_d_bfwt <= din_11_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_din_11_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_din_11_rsc_wait_ctrl
    (
  core_wen, core_wten, din_11_rsci_oswt, din_11_rsci_biwt, din_11_rsci_bdwt, din_11_rsci_biwt_pff,
      din_11_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_11_rsci_oswt;
  output din_11_rsci_biwt;
  output din_11_rsci_bdwt;
  output din_11_rsci_biwt_pff;
  input din_11_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_11_rsci_bdwt = din_11_rsci_oswt & core_wen;
  assign din_11_rsci_biwt = (~ core_wten) & din_11_rsci_oswt;
  assign din_11_rsci_biwt_pff = core_wen & din_11_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_din_10_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_din_10_rsc_wait_dp (
  clk, rst, din_10_rsci_douta_d, din_10_rsci_douta_d_mxwt, din_10_rsci_biwt, din_10_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_10_rsci_douta_d;
  output [63:0] din_10_rsci_douta_d_mxwt;
  input din_10_rsci_biwt;
  input din_10_rsci_bdwt;


  // Interconnect Declarations
  reg din_10_rsci_bcwt;
  reg [63:0] din_10_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_10_rsci_douta_d_mxwt = MUX_v_64_2_2(din_10_rsci_douta_d, din_10_rsci_douta_d_bfwt,
      din_10_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_10_rsci_bcwt <= 1'b0;
      din_10_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_10_rsci_bcwt <= ~((~(din_10_rsci_bcwt | din_10_rsci_biwt)) | din_10_rsci_bdwt);
      din_10_rsci_douta_d_bfwt <= din_10_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_din_10_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_din_10_rsc_wait_ctrl
    (
  core_wen, core_wten, din_10_rsci_oswt, din_10_rsci_biwt, din_10_rsci_bdwt, din_10_rsci_biwt_pff,
      din_10_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_10_rsci_oswt;
  output din_10_rsci_biwt;
  output din_10_rsci_bdwt;
  output din_10_rsci_biwt_pff;
  input din_10_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_10_rsci_bdwt = din_10_rsci_oswt & core_wen;
  assign din_10_rsci_biwt = (~ core_wten) & din_10_rsci_oswt;
  assign din_10_rsci_biwt_pff = core_wen & din_10_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_din_9_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_din_9_rsc_wait_dp (
  clk, rst, din_9_rsci_douta_d, din_9_rsci_douta_d_mxwt, din_9_rsci_biwt, din_9_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_9_rsci_douta_d;
  output [63:0] din_9_rsci_douta_d_mxwt;
  input din_9_rsci_biwt;
  input din_9_rsci_bdwt;


  // Interconnect Declarations
  reg din_9_rsci_bcwt;
  reg [63:0] din_9_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_9_rsci_douta_d_mxwt = MUX_v_64_2_2(din_9_rsci_douta_d, din_9_rsci_douta_d_bfwt,
      din_9_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_9_rsci_bcwt <= 1'b0;
      din_9_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_9_rsci_bcwt <= ~((~(din_9_rsci_bcwt | din_9_rsci_biwt)) | din_9_rsci_bdwt);
      din_9_rsci_douta_d_bfwt <= din_9_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_din_9_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_din_9_rsc_wait_ctrl (
  core_wen, core_wten, din_9_rsci_oswt, din_9_rsci_biwt, din_9_rsci_bdwt, din_9_rsci_biwt_pff,
      din_9_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_9_rsci_oswt;
  output din_9_rsci_biwt;
  output din_9_rsci_bdwt;
  output din_9_rsci_biwt_pff;
  input din_9_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_9_rsci_bdwt = din_9_rsci_oswt & core_wen;
  assign din_9_rsci_biwt = (~ core_wten) & din_9_rsci_oswt;
  assign din_9_rsci_biwt_pff = core_wen & din_9_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_din_8_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_din_8_rsc_wait_dp (
  clk, rst, din_8_rsci_douta_d, din_8_rsci_douta_d_mxwt, din_8_rsci_biwt, din_8_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_8_rsci_douta_d;
  output [63:0] din_8_rsci_douta_d_mxwt;
  input din_8_rsci_biwt;
  input din_8_rsci_bdwt;


  // Interconnect Declarations
  reg din_8_rsci_bcwt;
  reg [63:0] din_8_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_8_rsci_douta_d_mxwt = MUX_v_64_2_2(din_8_rsci_douta_d, din_8_rsci_douta_d_bfwt,
      din_8_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_8_rsci_bcwt <= 1'b0;
      din_8_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_8_rsci_bcwt <= ~((~(din_8_rsci_bcwt | din_8_rsci_biwt)) | din_8_rsci_bdwt);
      din_8_rsci_douta_d_bfwt <= din_8_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_din_8_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_din_8_rsc_wait_ctrl (
  core_wen, core_wten, din_8_rsci_oswt, din_8_rsci_biwt, din_8_rsci_bdwt, din_8_rsci_biwt_pff,
      din_8_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_8_rsci_oswt;
  output din_8_rsci_biwt;
  output din_8_rsci_bdwt;
  output din_8_rsci_biwt_pff;
  input din_8_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_8_rsci_bdwt = din_8_rsci_oswt & core_wen;
  assign din_8_rsci_biwt = (~ core_wten) & din_8_rsci_oswt;
  assign din_8_rsci_biwt_pff = core_wen & din_8_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_din_7_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_din_7_rsc_wait_dp (
  clk, rst, din_7_rsci_douta_d, din_7_rsci_douta_d_mxwt, din_7_rsci_biwt, din_7_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_7_rsci_douta_d;
  output [63:0] din_7_rsci_douta_d_mxwt;
  input din_7_rsci_biwt;
  input din_7_rsci_bdwt;


  // Interconnect Declarations
  reg din_7_rsci_bcwt;
  reg [63:0] din_7_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_7_rsci_douta_d_mxwt = MUX_v_64_2_2(din_7_rsci_douta_d, din_7_rsci_douta_d_bfwt,
      din_7_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_7_rsci_bcwt <= 1'b0;
      din_7_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_7_rsci_bcwt <= ~((~(din_7_rsci_bcwt | din_7_rsci_biwt)) | din_7_rsci_bdwt);
      din_7_rsci_douta_d_bfwt <= din_7_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_din_7_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_din_7_rsc_wait_ctrl (
  core_wen, core_wten, din_7_rsci_oswt, din_7_rsci_biwt, din_7_rsci_bdwt, din_7_rsci_biwt_pff,
      din_7_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_7_rsci_oswt;
  output din_7_rsci_biwt;
  output din_7_rsci_bdwt;
  output din_7_rsci_biwt_pff;
  input din_7_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_7_rsci_bdwt = din_7_rsci_oswt & core_wen;
  assign din_7_rsci_biwt = (~ core_wten) & din_7_rsci_oswt;
  assign din_7_rsci_biwt_pff = core_wen & din_7_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_din_6_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_din_6_rsc_wait_dp (
  clk, rst, din_6_rsci_douta_d, din_6_rsci_douta_d_mxwt, din_6_rsci_biwt, din_6_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_6_rsci_douta_d;
  output [63:0] din_6_rsci_douta_d_mxwt;
  input din_6_rsci_biwt;
  input din_6_rsci_bdwt;


  // Interconnect Declarations
  reg din_6_rsci_bcwt;
  reg [63:0] din_6_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_6_rsci_douta_d_mxwt = MUX_v_64_2_2(din_6_rsci_douta_d, din_6_rsci_douta_d_bfwt,
      din_6_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_6_rsci_bcwt <= 1'b0;
      din_6_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_6_rsci_bcwt <= ~((~(din_6_rsci_bcwt | din_6_rsci_biwt)) | din_6_rsci_bdwt);
      din_6_rsci_douta_d_bfwt <= din_6_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_din_6_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_din_6_rsc_wait_ctrl (
  core_wen, core_wten, din_6_rsci_oswt, din_6_rsci_biwt, din_6_rsci_bdwt, din_6_rsci_biwt_pff,
      din_6_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_6_rsci_oswt;
  output din_6_rsci_biwt;
  output din_6_rsci_bdwt;
  output din_6_rsci_biwt_pff;
  input din_6_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_6_rsci_bdwt = din_6_rsci_oswt & core_wen;
  assign din_6_rsci_biwt = (~ core_wten) & din_6_rsci_oswt;
  assign din_6_rsci_biwt_pff = core_wen & din_6_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_din_5_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_din_5_rsc_wait_dp (
  clk, rst, din_5_rsci_douta_d, din_5_rsci_douta_d_mxwt, din_5_rsci_biwt, din_5_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_5_rsci_douta_d;
  output [63:0] din_5_rsci_douta_d_mxwt;
  input din_5_rsci_biwt;
  input din_5_rsci_bdwt;


  // Interconnect Declarations
  reg din_5_rsci_bcwt;
  reg [63:0] din_5_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_5_rsci_douta_d_mxwt = MUX_v_64_2_2(din_5_rsci_douta_d, din_5_rsci_douta_d_bfwt,
      din_5_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_5_rsci_bcwt <= 1'b0;
      din_5_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_5_rsci_bcwt <= ~((~(din_5_rsci_bcwt | din_5_rsci_biwt)) | din_5_rsci_bdwt);
      din_5_rsci_douta_d_bfwt <= din_5_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_din_5_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_din_5_rsc_wait_ctrl (
  core_wen, core_wten, din_5_rsci_oswt, din_5_rsci_biwt, din_5_rsci_bdwt, din_5_rsci_biwt_pff,
      din_5_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_5_rsci_oswt;
  output din_5_rsci_biwt;
  output din_5_rsci_bdwt;
  output din_5_rsci_biwt_pff;
  input din_5_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_5_rsci_bdwt = din_5_rsci_oswt & core_wen;
  assign din_5_rsci_biwt = (~ core_wten) & din_5_rsci_oswt;
  assign din_5_rsci_biwt_pff = core_wen & din_5_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_din_4_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_din_4_rsc_wait_dp (
  clk, rst, din_4_rsci_douta_d, din_4_rsci_douta_d_mxwt, din_4_rsci_biwt, din_4_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_4_rsci_douta_d;
  output [63:0] din_4_rsci_douta_d_mxwt;
  input din_4_rsci_biwt;
  input din_4_rsci_bdwt;


  // Interconnect Declarations
  reg din_4_rsci_bcwt;
  reg [63:0] din_4_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_4_rsci_douta_d_mxwt = MUX_v_64_2_2(din_4_rsci_douta_d, din_4_rsci_douta_d_bfwt,
      din_4_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_4_rsci_bcwt <= 1'b0;
      din_4_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_4_rsci_bcwt <= ~((~(din_4_rsci_bcwt | din_4_rsci_biwt)) | din_4_rsci_bdwt);
      din_4_rsci_douta_d_bfwt <= din_4_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_din_4_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_din_4_rsc_wait_ctrl (
  core_wen, core_wten, din_4_rsci_oswt, din_4_rsci_biwt, din_4_rsci_bdwt, din_4_rsci_biwt_pff,
      din_4_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_4_rsci_oswt;
  output din_4_rsci_biwt;
  output din_4_rsci_bdwt;
  output din_4_rsci_biwt_pff;
  input din_4_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_4_rsci_bdwt = din_4_rsci_oswt & core_wen;
  assign din_4_rsci_biwt = (~ core_wten) & din_4_rsci_oswt;
  assign din_4_rsci_biwt_pff = core_wen & din_4_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_din_3_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_din_3_rsc_wait_dp (
  clk, rst, din_3_rsci_douta_d, din_3_rsci_douta_d_mxwt, din_3_rsci_biwt, din_3_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_3_rsci_douta_d;
  output [63:0] din_3_rsci_douta_d_mxwt;
  input din_3_rsci_biwt;
  input din_3_rsci_bdwt;


  // Interconnect Declarations
  reg din_3_rsci_bcwt;
  reg [63:0] din_3_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_3_rsci_douta_d_mxwt = MUX_v_64_2_2(din_3_rsci_douta_d, din_3_rsci_douta_d_bfwt,
      din_3_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_3_rsci_bcwt <= 1'b0;
      din_3_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_3_rsci_bcwt <= ~((~(din_3_rsci_bcwt | din_3_rsci_biwt)) | din_3_rsci_bdwt);
      din_3_rsci_douta_d_bfwt <= din_3_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_din_3_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_din_3_rsc_wait_ctrl (
  core_wen, core_wten, din_3_rsci_oswt, din_3_rsci_biwt, din_3_rsci_bdwt, din_3_rsci_biwt_pff,
      din_3_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_3_rsci_oswt;
  output din_3_rsci_biwt;
  output din_3_rsci_bdwt;
  output din_3_rsci_biwt_pff;
  input din_3_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_3_rsci_bdwt = din_3_rsci_oswt & core_wen;
  assign din_3_rsci_biwt = (~ core_wten) & din_3_rsci_oswt;
  assign din_3_rsci_biwt_pff = core_wen & din_3_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_din_2_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_din_2_rsc_wait_dp (
  clk, rst, din_2_rsci_douta_d, din_2_rsci_douta_d_mxwt, din_2_rsci_biwt, din_2_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_2_rsci_douta_d;
  output [63:0] din_2_rsci_douta_d_mxwt;
  input din_2_rsci_biwt;
  input din_2_rsci_bdwt;


  // Interconnect Declarations
  reg din_2_rsci_bcwt;
  reg [63:0] din_2_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_2_rsci_douta_d_mxwt = MUX_v_64_2_2(din_2_rsci_douta_d, din_2_rsci_douta_d_bfwt,
      din_2_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_2_rsci_bcwt <= 1'b0;
      din_2_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_2_rsci_bcwt <= ~((~(din_2_rsci_bcwt | din_2_rsci_biwt)) | din_2_rsci_bdwt);
      din_2_rsci_douta_d_bfwt <= din_2_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_din_2_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_din_2_rsc_wait_ctrl (
  core_wen, core_wten, din_2_rsci_oswt, din_2_rsci_biwt, din_2_rsci_bdwt, din_2_rsci_biwt_pff,
      din_2_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_2_rsci_oswt;
  output din_2_rsci_biwt;
  output din_2_rsci_bdwt;
  output din_2_rsci_biwt_pff;
  input din_2_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_2_rsci_bdwt = din_2_rsci_oswt & core_wen;
  assign din_2_rsci_biwt = (~ core_wten) & din_2_rsci_oswt;
  assign din_2_rsci_biwt_pff = core_wen & din_2_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_din_1_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_din_1_rsc_wait_dp (
  clk, rst, din_1_rsci_douta_d, din_1_rsci_douta_d_mxwt, din_1_rsci_biwt, din_1_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_1_rsci_douta_d;
  output [63:0] din_1_rsci_douta_d_mxwt;
  input din_1_rsci_biwt;
  input din_1_rsci_bdwt;


  // Interconnect Declarations
  reg din_1_rsci_bcwt;
  reg [63:0] din_1_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_1_rsci_douta_d_mxwt = MUX_v_64_2_2(din_1_rsci_douta_d, din_1_rsci_douta_d_bfwt,
      din_1_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_1_rsci_bcwt <= 1'b0;
      din_1_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_1_rsci_bcwt <= ~((~(din_1_rsci_bcwt | din_1_rsci_biwt)) | din_1_rsci_bdwt);
      din_1_rsci_douta_d_bfwt <= din_1_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_din_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_din_1_rsc_wait_ctrl (
  core_wen, core_wten, din_1_rsci_oswt, din_1_rsci_biwt, din_1_rsci_bdwt, din_1_rsci_biwt_pff,
      din_1_rsci_oswt_pff
);
  input core_wen;
  input core_wten;
  input din_1_rsci_oswt;
  output din_1_rsci_biwt;
  output din_1_rsci_bdwt;
  output din_1_rsci_biwt_pff;
  input din_1_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_1_rsci_bdwt = din_1_rsci_oswt & core_wen;
  assign din_1_rsci_biwt = (~ core_wten) & din_1_rsci_oswt;
  assign din_1_rsci_biwt_pff = core_wen & din_1_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_din_0_rsc_wait_dp
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_din_0_rsc_wait_dp (
  clk, rst, din_0_rsci_douta_d, din_0_rsci_douta_d_mxwt, din_0_rsci_biwt, din_0_rsci_bdwt
);
  input clk;
  input rst;
  input [63:0] din_0_rsci_douta_d;
  output [63:0] din_0_rsci_douta_d_mxwt;
  input din_0_rsci_biwt;
  input din_0_rsci_bdwt;


  // Interconnect Declarations
  reg din_0_rsci_bcwt;
  reg [63:0] din_0_rsci_douta_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_0_rsci_douta_d_mxwt = MUX_v_64_2_2(din_0_rsci_douta_d, din_0_rsci_douta_d_bfwt,
      din_0_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      din_0_rsci_bcwt <= 1'b0;
      din_0_rsci_douta_d_bfwt <= 64'b0;
    end
    else begin
      din_0_rsci_bcwt <= ~((~(din_0_rsci_bcwt | din_0_rsci_biwt)) | din_0_rsci_bdwt);
      din_0_rsci_douta_d_bfwt <= din_0_rsci_douta_d_mxwt;
    end
  end

  function [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_din_0_rsc_wait_ctrl
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_din_0_rsc_wait_ctrl (
  core_wen, din_0_rsci_oswt, core_wten, din_0_rsci_biwt, din_0_rsci_bdwt, din_0_rsci_biwt_pff,
      din_0_rsci_oswt_pff
);
  input core_wen;
  input din_0_rsci_oswt;
  input core_wten;
  output din_0_rsci_biwt;
  output din_0_rsci_bdwt;
  output din_0_rsci_biwt_pff;
  input din_0_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_0_rsci_bdwt = din_0_rsci_oswt & core_wen;
  assign din_0_rsci_biwt = (~ core_wten) & din_0_rsci_oswt;
  assign din_0_rsci_biwt_pff = core_wen & din_0_rsci_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj (
  clk, rst, dout_0_rsc_req_vz, core_wen, core_wten, dout_0_rsc_req_obj_oswt, dout_0_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_0_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_0_rsc_req_obj_oswt;
  output dout_0_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_0_rsc_req_obj_vd;
  wire dout_0_rsc_req_obj_biwt;
  wire dout_0_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_0_rsc_req_obj (
      .vd(dout_0_rsc_req_obj_vd),
      .vz(dout_0_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_0_rsc_req_obj_oswt(dout_0_rsc_req_obj_oswt),
      .dout_0_rsc_req_obj_vd(dout_0_rsc_req_obj_vd),
      .dout_0_rsc_req_obj_biwt(dout_0_rsc_req_obj_biwt),
      .dout_0_rsc_req_obj_bdwt(dout_0_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_0_rsc_req_obj_oswt(dout_0_rsc_req_obj_oswt),
      .dout_0_rsc_req_obj_wen_comp(dout_0_rsc_req_obj_wen_comp),
      .dout_0_rsc_req_obj_biwt(dout_0_rsc_req_obj_biwt),
      .dout_0_rsc_req_obj_bdwt(dout_0_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_rls_obj (
  dout_0_rsc_rls_lz, core_wten, dout_0_rsc_rls_obj_iswt0
);
  output dout_0_rsc_rls_lz;
  input core_wten;
  input dout_0_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_0_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_0_rsc_rls_obj (
      .ld(dout_0_rsc_rls_obj_ld_core_sct),
      .lz(dout_0_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_rls_obj_dout_0_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_rls_obj_dout_0_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_0_rsc_rls_obj_iswt0(dout_0_rsc_rls_obj_iswt0),
      .dout_0_rsc_rls_obj_ld_core_sct(dout_0_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj (
  clk, rst, dout_1_rsc_req_vz, core_wen, core_wten, dout_1_rsc_req_obj_oswt, dout_1_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_1_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_1_rsc_req_obj_oswt;
  output dout_1_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_1_rsc_req_obj_vd;
  wire dout_1_rsc_req_obj_biwt;
  wire dout_1_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_1_rsc_req_obj (
      .vd(dout_1_rsc_req_obj_vd),
      .vz(dout_1_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_1_rsc_req_obj_oswt(dout_1_rsc_req_obj_oswt),
      .dout_1_rsc_req_obj_vd(dout_1_rsc_req_obj_vd),
      .dout_1_rsc_req_obj_biwt(dout_1_rsc_req_obj_biwt),
      .dout_1_rsc_req_obj_bdwt(dout_1_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_1_rsc_req_obj_oswt(dout_1_rsc_req_obj_oswt),
      .dout_1_rsc_req_obj_wen_comp(dout_1_rsc_req_obj_wen_comp),
      .dout_1_rsc_req_obj_biwt(dout_1_rsc_req_obj_biwt),
      .dout_1_rsc_req_obj_bdwt(dout_1_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_rls_obj (
  dout_1_rsc_rls_lz, core_wten, dout_1_rsc_rls_obj_iswt0
);
  output dout_1_rsc_rls_lz;
  input core_wten;
  input dout_1_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_1_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_1_rsc_rls_obj (
      .ld(dout_1_rsc_rls_obj_ld_core_sct),
      .lz(dout_1_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_rls_obj_dout_1_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_rls_obj_dout_1_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_1_rsc_rls_obj_iswt0(dout_1_rsc_rls_obj_iswt0),
      .dout_1_rsc_rls_obj_ld_core_sct(dout_1_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj (
  clk, rst, dout_2_rsc_req_vz, core_wen, core_wten, dout_2_rsc_req_obj_oswt, dout_2_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_2_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_2_rsc_req_obj_oswt;
  output dout_2_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_2_rsc_req_obj_vd;
  wire dout_2_rsc_req_obj_biwt;
  wire dout_2_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_2_rsc_req_obj (
      .vd(dout_2_rsc_req_obj_vd),
      .vz(dout_2_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_2_rsc_req_obj_oswt(dout_2_rsc_req_obj_oswt),
      .dout_2_rsc_req_obj_vd(dout_2_rsc_req_obj_vd),
      .dout_2_rsc_req_obj_biwt(dout_2_rsc_req_obj_biwt),
      .dout_2_rsc_req_obj_bdwt(dout_2_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_2_rsc_req_obj_oswt(dout_2_rsc_req_obj_oswt),
      .dout_2_rsc_req_obj_wen_comp(dout_2_rsc_req_obj_wen_comp),
      .dout_2_rsc_req_obj_biwt(dout_2_rsc_req_obj_biwt),
      .dout_2_rsc_req_obj_bdwt(dout_2_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_rls_obj (
  dout_2_rsc_rls_lz, core_wten, dout_2_rsc_rls_obj_iswt0
);
  output dout_2_rsc_rls_lz;
  input core_wten;
  input dout_2_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_2_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_2_rsc_rls_obj (
      .ld(dout_2_rsc_rls_obj_ld_core_sct),
      .lz(dout_2_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_rls_obj_dout_2_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_rls_obj_dout_2_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_2_rsc_rls_obj_iswt0(dout_2_rsc_rls_obj_iswt0),
      .dout_2_rsc_rls_obj_ld_core_sct(dout_2_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj (
  clk, rst, dout_3_rsc_req_vz, core_wen, core_wten, dout_3_rsc_req_obj_oswt, dout_3_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_3_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_3_rsc_req_obj_oswt;
  output dout_3_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_3_rsc_req_obj_vd;
  wire dout_3_rsc_req_obj_biwt;
  wire dout_3_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_3_rsc_req_obj (
      .vd(dout_3_rsc_req_obj_vd),
      .vz(dout_3_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_3_rsc_req_obj_oswt(dout_3_rsc_req_obj_oswt),
      .dout_3_rsc_req_obj_vd(dout_3_rsc_req_obj_vd),
      .dout_3_rsc_req_obj_biwt(dout_3_rsc_req_obj_biwt),
      .dout_3_rsc_req_obj_bdwt(dout_3_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_3_rsc_req_obj_oswt(dout_3_rsc_req_obj_oswt),
      .dout_3_rsc_req_obj_wen_comp(dout_3_rsc_req_obj_wen_comp),
      .dout_3_rsc_req_obj_biwt(dout_3_rsc_req_obj_biwt),
      .dout_3_rsc_req_obj_bdwt(dout_3_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_rls_obj (
  dout_3_rsc_rls_lz, core_wten, dout_3_rsc_rls_obj_iswt0
);
  output dout_3_rsc_rls_lz;
  input core_wten;
  input dout_3_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_3_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_3_rsc_rls_obj (
      .ld(dout_3_rsc_rls_obj_ld_core_sct),
      .lz(dout_3_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_rls_obj_dout_3_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_rls_obj_dout_3_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_3_rsc_rls_obj_iswt0(dout_3_rsc_rls_obj_iswt0),
      .dout_3_rsc_rls_obj_ld_core_sct(dout_3_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj (
  clk, rst, dout_4_rsc_req_vz, core_wen, core_wten, dout_4_rsc_req_obj_oswt, dout_4_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_4_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_4_rsc_req_obj_oswt;
  output dout_4_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_4_rsc_req_obj_vd;
  wire dout_4_rsc_req_obj_biwt;
  wire dout_4_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_4_rsc_req_obj (
      .vd(dout_4_rsc_req_obj_vd),
      .vz(dout_4_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_4_rsc_req_obj_oswt(dout_4_rsc_req_obj_oswt),
      .dout_4_rsc_req_obj_vd(dout_4_rsc_req_obj_vd),
      .dout_4_rsc_req_obj_biwt(dout_4_rsc_req_obj_biwt),
      .dout_4_rsc_req_obj_bdwt(dout_4_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_4_rsc_req_obj_oswt(dout_4_rsc_req_obj_oswt),
      .dout_4_rsc_req_obj_wen_comp(dout_4_rsc_req_obj_wen_comp),
      .dout_4_rsc_req_obj_biwt(dout_4_rsc_req_obj_biwt),
      .dout_4_rsc_req_obj_bdwt(dout_4_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_rls_obj (
  dout_4_rsc_rls_lz, core_wten, dout_4_rsc_rls_obj_iswt0
);
  output dout_4_rsc_rls_lz;
  input core_wten;
  input dout_4_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_4_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_4_rsc_rls_obj (
      .ld(dout_4_rsc_rls_obj_ld_core_sct),
      .lz(dout_4_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_rls_obj_dout_4_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_rls_obj_dout_4_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_4_rsc_rls_obj_iswt0(dout_4_rsc_rls_obj_iswt0),
      .dout_4_rsc_rls_obj_ld_core_sct(dout_4_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj (
  clk, rst, dout_5_rsc_req_vz, core_wen, core_wten, dout_5_rsc_req_obj_oswt, dout_5_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_5_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_5_rsc_req_obj_oswt;
  output dout_5_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_5_rsc_req_obj_vd;
  wire dout_5_rsc_req_obj_biwt;
  wire dout_5_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_5_rsc_req_obj (
      .vd(dout_5_rsc_req_obj_vd),
      .vz(dout_5_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_5_rsc_req_obj_oswt(dout_5_rsc_req_obj_oswt),
      .dout_5_rsc_req_obj_vd(dout_5_rsc_req_obj_vd),
      .dout_5_rsc_req_obj_biwt(dout_5_rsc_req_obj_biwt),
      .dout_5_rsc_req_obj_bdwt(dout_5_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_5_rsc_req_obj_oswt(dout_5_rsc_req_obj_oswt),
      .dout_5_rsc_req_obj_wen_comp(dout_5_rsc_req_obj_wen_comp),
      .dout_5_rsc_req_obj_biwt(dout_5_rsc_req_obj_biwt),
      .dout_5_rsc_req_obj_bdwt(dout_5_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_rls_obj (
  dout_5_rsc_rls_lz, core_wten, dout_5_rsc_rls_obj_iswt0
);
  output dout_5_rsc_rls_lz;
  input core_wten;
  input dout_5_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_5_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_5_rsc_rls_obj (
      .ld(dout_5_rsc_rls_obj_ld_core_sct),
      .lz(dout_5_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_rls_obj_dout_5_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_rls_obj_dout_5_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_5_rsc_rls_obj_iswt0(dout_5_rsc_rls_obj_iswt0),
      .dout_5_rsc_rls_obj_ld_core_sct(dout_5_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj (
  clk, rst, dout_6_rsc_req_vz, core_wen, core_wten, dout_6_rsc_req_obj_oswt, dout_6_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_6_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_6_rsc_req_obj_oswt;
  output dout_6_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_6_rsc_req_obj_vd;
  wire dout_6_rsc_req_obj_biwt;
  wire dout_6_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_6_rsc_req_obj (
      .vd(dout_6_rsc_req_obj_vd),
      .vz(dout_6_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_6_rsc_req_obj_oswt(dout_6_rsc_req_obj_oswt),
      .dout_6_rsc_req_obj_vd(dout_6_rsc_req_obj_vd),
      .dout_6_rsc_req_obj_biwt(dout_6_rsc_req_obj_biwt),
      .dout_6_rsc_req_obj_bdwt(dout_6_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_6_rsc_req_obj_oswt(dout_6_rsc_req_obj_oswt),
      .dout_6_rsc_req_obj_wen_comp(dout_6_rsc_req_obj_wen_comp),
      .dout_6_rsc_req_obj_biwt(dout_6_rsc_req_obj_biwt),
      .dout_6_rsc_req_obj_bdwt(dout_6_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_rls_obj (
  dout_6_rsc_rls_lz, core_wten, dout_6_rsc_rls_obj_iswt0
);
  output dout_6_rsc_rls_lz;
  input core_wten;
  input dout_6_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_6_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_6_rsc_rls_obj (
      .ld(dout_6_rsc_rls_obj_ld_core_sct),
      .lz(dout_6_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_rls_obj_dout_6_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_rls_obj_dout_6_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_6_rsc_rls_obj_iswt0(dout_6_rsc_rls_obj_iswt0),
      .dout_6_rsc_rls_obj_ld_core_sct(dout_6_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj (
  clk, rst, dout_7_rsc_req_vz, core_wen, core_wten, dout_7_rsc_req_obj_oswt, dout_7_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_7_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_7_rsc_req_obj_oswt;
  output dout_7_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_7_rsc_req_obj_vd;
  wire dout_7_rsc_req_obj_biwt;
  wire dout_7_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_7_rsc_req_obj (
      .vd(dout_7_rsc_req_obj_vd),
      .vz(dout_7_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_7_rsc_req_obj_oswt(dout_7_rsc_req_obj_oswt),
      .dout_7_rsc_req_obj_vd(dout_7_rsc_req_obj_vd),
      .dout_7_rsc_req_obj_biwt(dout_7_rsc_req_obj_biwt),
      .dout_7_rsc_req_obj_bdwt(dout_7_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_7_rsc_req_obj_oswt(dout_7_rsc_req_obj_oswt),
      .dout_7_rsc_req_obj_wen_comp(dout_7_rsc_req_obj_wen_comp),
      .dout_7_rsc_req_obj_biwt(dout_7_rsc_req_obj_biwt),
      .dout_7_rsc_req_obj_bdwt(dout_7_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_rls_obj (
  dout_7_rsc_rls_lz, core_wten, dout_7_rsc_rls_obj_iswt0
);
  output dout_7_rsc_rls_lz;
  input core_wten;
  input dout_7_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_7_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_7_rsc_rls_obj (
      .ld(dout_7_rsc_rls_obj_ld_core_sct),
      .lz(dout_7_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_rls_obj_dout_7_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_rls_obj_dout_7_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_7_rsc_rls_obj_iswt0(dout_7_rsc_rls_obj_iswt0),
      .dout_7_rsc_rls_obj_ld_core_sct(dout_7_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj (
  clk, rst, dout_8_rsc_req_vz, core_wen, core_wten, dout_8_rsc_req_obj_oswt, dout_8_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_8_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_8_rsc_req_obj_oswt;
  output dout_8_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_8_rsc_req_obj_vd;
  wire dout_8_rsc_req_obj_biwt;
  wire dout_8_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_8_rsc_req_obj (
      .vd(dout_8_rsc_req_obj_vd),
      .vz(dout_8_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_8_rsc_req_obj_oswt(dout_8_rsc_req_obj_oswt),
      .dout_8_rsc_req_obj_vd(dout_8_rsc_req_obj_vd),
      .dout_8_rsc_req_obj_biwt(dout_8_rsc_req_obj_biwt),
      .dout_8_rsc_req_obj_bdwt(dout_8_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_8_rsc_req_obj_oswt(dout_8_rsc_req_obj_oswt),
      .dout_8_rsc_req_obj_wen_comp(dout_8_rsc_req_obj_wen_comp),
      .dout_8_rsc_req_obj_biwt(dout_8_rsc_req_obj_biwt),
      .dout_8_rsc_req_obj_bdwt(dout_8_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_rls_obj (
  dout_8_rsc_rls_lz, core_wten, dout_8_rsc_rls_obj_iswt0
);
  output dout_8_rsc_rls_lz;
  input core_wten;
  input dout_8_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_8_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_8_rsc_rls_obj (
      .ld(dout_8_rsc_rls_obj_ld_core_sct),
      .lz(dout_8_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_rls_obj_dout_8_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_rls_obj_dout_8_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_8_rsc_rls_obj_iswt0(dout_8_rsc_rls_obj_iswt0),
      .dout_8_rsc_rls_obj_ld_core_sct(dout_8_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj (
  clk, rst, dout_9_rsc_req_vz, core_wen, core_wten, dout_9_rsc_req_obj_oswt, dout_9_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_9_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_9_rsc_req_obj_oswt;
  output dout_9_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_9_rsc_req_obj_vd;
  wire dout_9_rsc_req_obj_biwt;
  wire dout_9_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_9_rsc_req_obj (
      .vd(dout_9_rsc_req_obj_vd),
      .vz(dout_9_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_9_rsc_req_obj_oswt(dout_9_rsc_req_obj_oswt),
      .dout_9_rsc_req_obj_vd(dout_9_rsc_req_obj_vd),
      .dout_9_rsc_req_obj_biwt(dout_9_rsc_req_obj_biwt),
      .dout_9_rsc_req_obj_bdwt(dout_9_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_9_rsc_req_obj_oswt(dout_9_rsc_req_obj_oswt),
      .dout_9_rsc_req_obj_wen_comp(dout_9_rsc_req_obj_wen_comp),
      .dout_9_rsc_req_obj_biwt(dout_9_rsc_req_obj_biwt),
      .dout_9_rsc_req_obj_bdwt(dout_9_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_rls_obj (
  dout_9_rsc_rls_lz, core_wten, dout_9_rsc_rls_obj_iswt0
);
  output dout_9_rsc_rls_lz;
  input core_wten;
  input dout_9_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_9_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_9_rsc_rls_obj (
      .ld(dout_9_rsc_rls_obj_ld_core_sct),
      .lz(dout_9_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_rls_obj_dout_9_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_rls_obj_dout_9_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_9_rsc_rls_obj_iswt0(dout_9_rsc_rls_obj_iswt0),
      .dout_9_rsc_rls_obj_ld_core_sct(dout_9_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj (
  clk, rst, dout_10_rsc_req_vz, core_wen, core_wten, dout_10_rsc_req_obj_oswt, dout_10_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_10_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_10_rsc_req_obj_oswt;
  output dout_10_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_10_rsc_req_obj_vd;
  wire dout_10_rsc_req_obj_biwt;
  wire dout_10_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_10_rsc_req_obj (
      .vd(dout_10_rsc_req_obj_vd),
      .vz(dout_10_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_10_rsc_req_obj_oswt(dout_10_rsc_req_obj_oswt),
      .dout_10_rsc_req_obj_vd(dout_10_rsc_req_obj_vd),
      .dout_10_rsc_req_obj_biwt(dout_10_rsc_req_obj_biwt),
      .dout_10_rsc_req_obj_bdwt(dout_10_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_10_rsc_req_obj_oswt(dout_10_rsc_req_obj_oswt),
      .dout_10_rsc_req_obj_wen_comp(dout_10_rsc_req_obj_wen_comp),
      .dout_10_rsc_req_obj_biwt(dout_10_rsc_req_obj_biwt),
      .dout_10_rsc_req_obj_bdwt(dout_10_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_rls_obj (
  dout_10_rsc_rls_lz, core_wten, dout_10_rsc_rls_obj_iswt0
);
  output dout_10_rsc_rls_lz;
  input core_wten;
  input dout_10_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_10_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_10_rsc_rls_obj (
      .ld(dout_10_rsc_rls_obj_ld_core_sct),
      .lz(dout_10_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_rls_obj_dout_10_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_rls_obj_dout_10_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_10_rsc_rls_obj_iswt0(dout_10_rsc_rls_obj_iswt0),
      .dout_10_rsc_rls_obj_ld_core_sct(dout_10_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj (
  clk, rst, dout_11_rsc_req_vz, core_wen, core_wten, dout_11_rsc_req_obj_oswt, dout_11_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_11_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_11_rsc_req_obj_oswt;
  output dout_11_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_11_rsc_req_obj_vd;
  wire dout_11_rsc_req_obj_biwt;
  wire dout_11_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_11_rsc_req_obj (
      .vd(dout_11_rsc_req_obj_vd),
      .vz(dout_11_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_11_rsc_req_obj_oswt(dout_11_rsc_req_obj_oswt),
      .dout_11_rsc_req_obj_vd(dout_11_rsc_req_obj_vd),
      .dout_11_rsc_req_obj_biwt(dout_11_rsc_req_obj_biwt),
      .dout_11_rsc_req_obj_bdwt(dout_11_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_11_rsc_req_obj_oswt(dout_11_rsc_req_obj_oswt),
      .dout_11_rsc_req_obj_wen_comp(dout_11_rsc_req_obj_wen_comp),
      .dout_11_rsc_req_obj_biwt(dout_11_rsc_req_obj_biwt),
      .dout_11_rsc_req_obj_bdwt(dout_11_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_rls_obj (
  dout_11_rsc_rls_lz, core_wten, dout_11_rsc_rls_obj_iswt0
);
  output dout_11_rsc_rls_lz;
  input core_wten;
  input dout_11_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_11_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_11_rsc_rls_obj (
      .ld(dout_11_rsc_rls_obj_ld_core_sct),
      .lz(dout_11_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_rls_obj_dout_11_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_rls_obj_dout_11_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_11_rsc_rls_obj_iswt0(dout_11_rsc_rls_obj_iswt0),
      .dout_11_rsc_rls_obj_ld_core_sct(dout_11_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj (
  clk, rst, dout_12_rsc_req_vz, core_wen, core_wten, dout_12_rsc_req_obj_oswt, dout_12_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_12_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_12_rsc_req_obj_oswt;
  output dout_12_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_12_rsc_req_obj_vd;
  wire dout_12_rsc_req_obj_biwt;
  wire dout_12_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_12_rsc_req_obj (
      .vd(dout_12_rsc_req_obj_vd),
      .vz(dout_12_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_12_rsc_req_obj_oswt(dout_12_rsc_req_obj_oswt),
      .dout_12_rsc_req_obj_vd(dout_12_rsc_req_obj_vd),
      .dout_12_rsc_req_obj_biwt(dout_12_rsc_req_obj_biwt),
      .dout_12_rsc_req_obj_bdwt(dout_12_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_12_rsc_req_obj_oswt(dout_12_rsc_req_obj_oswt),
      .dout_12_rsc_req_obj_wen_comp(dout_12_rsc_req_obj_wen_comp),
      .dout_12_rsc_req_obj_biwt(dout_12_rsc_req_obj_biwt),
      .dout_12_rsc_req_obj_bdwt(dout_12_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_rls_obj (
  dout_12_rsc_rls_lz, core_wten, dout_12_rsc_rls_obj_iswt0
);
  output dout_12_rsc_rls_lz;
  input core_wten;
  input dout_12_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_12_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_12_rsc_rls_obj (
      .ld(dout_12_rsc_rls_obj_ld_core_sct),
      .lz(dout_12_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_rls_obj_dout_12_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_rls_obj_dout_12_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_12_rsc_rls_obj_iswt0(dout_12_rsc_rls_obj_iswt0),
      .dout_12_rsc_rls_obj_ld_core_sct(dout_12_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj (
  clk, rst, dout_13_rsc_req_vz, core_wen, core_wten, dout_13_rsc_req_obj_oswt, dout_13_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_13_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_13_rsc_req_obj_oswt;
  output dout_13_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_13_rsc_req_obj_vd;
  wire dout_13_rsc_req_obj_biwt;
  wire dout_13_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_13_rsc_req_obj (
      .vd(dout_13_rsc_req_obj_vd),
      .vz(dout_13_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_13_rsc_req_obj_oswt(dout_13_rsc_req_obj_oswt),
      .dout_13_rsc_req_obj_vd(dout_13_rsc_req_obj_vd),
      .dout_13_rsc_req_obj_biwt(dout_13_rsc_req_obj_biwt),
      .dout_13_rsc_req_obj_bdwt(dout_13_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_13_rsc_req_obj_oswt(dout_13_rsc_req_obj_oswt),
      .dout_13_rsc_req_obj_wen_comp(dout_13_rsc_req_obj_wen_comp),
      .dout_13_rsc_req_obj_biwt(dout_13_rsc_req_obj_biwt),
      .dout_13_rsc_req_obj_bdwt(dout_13_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_rls_obj (
  dout_13_rsc_rls_lz, core_wten, dout_13_rsc_rls_obj_iswt0
);
  output dout_13_rsc_rls_lz;
  input core_wten;
  input dout_13_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_13_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_13_rsc_rls_obj (
      .ld(dout_13_rsc_rls_obj_ld_core_sct),
      .lz(dout_13_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_rls_obj_dout_13_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_rls_obj_dout_13_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_13_rsc_rls_obj_iswt0(dout_13_rsc_rls_obj_iswt0),
      .dout_13_rsc_rls_obj_ld_core_sct(dout_13_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj (
  clk, rst, dout_14_rsc_req_vz, core_wen, core_wten, dout_14_rsc_req_obj_oswt, dout_14_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_14_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_14_rsc_req_obj_oswt;
  output dout_14_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_14_rsc_req_obj_vd;
  wire dout_14_rsc_req_obj_biwt;
  wire dout_14_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_14_rsc_req_obj (
      .vd(dout_14_rsc_req_obj_vd),
      .vz(dout_14_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_14_rsc_req_obj_oswt(dout_14_rsc_req_obj_oswt),
      .dout_14_rsc_req_obj_vd(dout_14_rsc_req_obj_vd),
      .dout_14_rsc_req_obj_biwt(dout_14_rsc_req_obj_biwt),
      .dout_14_rsc_req_obj_bdwt(dout_14_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_14_rsc_req_obj_oswt(dout_14_rsc_req_obj_oswt),
      .dout_14_rsc_req_obj_wen_comp(dout_14_rsc_req_obj_wen_comp),
      .dout_14_rsc_req_obj_biwt(dout_14_rsc_req_obj_biwt),
      .dout_14_rsc_req_obj_bdwt(dout_14_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_rls_obj (
  dout_14_rsc_rls_lz, core_wten, dout_14_rsc_rls_obj_iswt0
);
  output dout_14_rsc_rls_lz;
  input core_wten;
  input dout_14_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_14_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_14_rsc_rls_obj (
      .ld(dout_14_rsc_rls_obj_ld_core_sct),
      .lz(dout_14_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_rls_obj_dout_14_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_rls_obj_dout_14_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_14_rsc_rls_obj_iswt0(dout_14_rsc_rls_obj_iswt0),
      .dout_14_rsc_rls_obj_ld_core_sct(dout_14_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj (
  clk, rst, dout_15_rsc_req_vz, core_wen, core_wten, dout_15_rsc_req_obj_oswt, dout_15_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_15_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_15_rsc_req_obj_oswt;
  output dout_15_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_15_rsc_req_obj_vd;
  wire dout_15_rsc_req_obj_biwt;
  wire dout_15_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_15_rsc_req_obj (
      .vd(dout_15_rsc_req_obj_vd),
      .vz(dout_15_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_15_rsc_req_obj_oswt(dout_15_rsc_req_obj_oswt),
      .dout_15_rsc_req_obj_vd(dout_15_rsc_req_obj_vd),
      .dout_15_rsc_req_obj_biwt(dout_15_rsc_req_obj_biwt),
      .dout_15_rsc_req_obj_bdwt(dout_15_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_15_rsc_req_obj_oswt(dout_15_rsc_req_obj_oswt),
      .dout_15_rsc_req_obj_wen_comp(dout_15_rsc_req_obj_wen_comp),
      .dout_15_rsc_req_obj_biwt(dout_15_rsc_req_obj_biwt),
      .dout_15_rsc_req_obj_bdwt(dout_15_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_rls_obj (
  dout_15_rsc_rls_lz, core_wten, dout_15_rsc_rls_obj_iswt0
);
  output dout_15_rsc_rls_lz;
  input core_wten;
  input dout_15_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_15_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_15_rsc_rls_obj (
      .ld(dout_15_rsc_rls_obj_ld_core_sct),
      .lz(dout_15_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_rls_obj_dout_15_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_rls_obj_dout_15_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_15_rsc_rls_obj_iswt0(dout_15_rsc_rls_obj_iswt0),
      .dout_15_rsc_rls_obj_ld_core_sct(dout_15_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj (
  clk, rst, dout_16_rsc_req_vz, core_wen, core_wten, dout_16_rsc_req_obj_oswt, dout_16_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_16_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_16_rsc_req_obj_oswt;
  output dout_16_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_16_rsc_req_obj_vd;
  wire dout_16_rsc_req_obj_biwt;
  wire dout_16_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_16_rsc_req_obj (
      .vd(dout_16_rsc_req_obj_vd),
      .vz(dout_16_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj_dout_16_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj_dout_16_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_16_rsc_req_obj_oswt(dout_16_rsc_req_obj_oswt),
      .dout_16_rsc_req_obj_vd(dout_16_rsc_req_obj_vd),
      .dout_16_rsc_req_obj_biwt(dout_16_rsc_req_obj_biwt),
      .dout_16_rsc_req_obj_bdwt(dout_16_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj_dout_16_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj_dout_16_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_16_rsc_req_obj_oswt(dout_16_rsc_req_obj_oswt),
      .dout_16_rsc_req_obj_wen_comp(dout_16_rsc_req_obj_wen_comp),
      .dout_16_rsc_req_obj_biwt(dout_16_rsc_req_obj_biwt),
      .dout_16_rsc_req_obj_bdwt(dout_16_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_rls_obj (
  dout_16_rsc_rls_lz, core_wten, dout_16_rsc_rls_obj_iswt0
);
  output dout_16_rsc_rls_lz;
  input core_wten;
  input dout_16_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_16_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_16_rsc_rls_obj (
      .ld(dout_16_rsc_rls_obj_ld_core_sct),
      .lz(dout_16_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_rls_obj_dout_16_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_rls_obj_dout_16_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_16_rsc_rls_obj_iswt0(dout_16_rsc_rls_obj_iswt0),
      .dout_16_rsc_rls_obj_ld_core_sct(dout_16_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj (
  clk, rst, dout_17_rsc_req_vz, core_wen, core_wten, dout_17_rsc_req_obj_oswt, dout_17_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_17_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_17_rsc_req_obj_oswt;
  output dout_17_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_17_rsc_req_obj_vd;
  wire dout_17_rsc_req_obj_biwt;
  wire dout_17_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_17_rsc_req_obj (
      .vd(dout_17_rsc_req_obj_vd),
      .vz(dout_17_rsc_req_vz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj_dout_17_rsc_req_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj_dout_17_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_17_rsc_req_obj_oswt(dout_17_rsc_req_obj_oswt),
      .dout_17_rsc_req_obj_vd(dout_17_rsc_req_obj_vd),
      .dout_17_rsc_req_obj_biwt(dout_17_rsc_req_obj_biwt),
      .dout_17_rsc_req_obj_bdwt(dout_17_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj_dout_17_rsc_req_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj_dout_17_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_17_rsc_req_obj_oswt(dout_17_rsc_req_obj_oswt),
      .dout_17_rsc_req_obj_wen_comp(dout_17_rsc_req_obj_wen_comp),
      .dout_17_rsc_req_obj_biwt(dout_17_rsc_req_obj_biwt),
      .dout_17_rsc_req_obj_bdwt(dout_17_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_rls_obj (
  dout_17_rsc_rls_lz, core_wten, dout_17_rsc_rls_obj_iswt0
);
  output dout_17_rsc_rls_lz;
  input core_wten;
  input dout_17_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_17_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_17_rsc_rls_obj (
      .ld(dout_17_rsc_rls_obj_ld_core_sct),
      .lz(dout_17_rsc_rls_lz)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_rls_obj_dout_17_rsc_rls_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_rls_obj_dout_17_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_17_rsc_rls_obj_iswt0(dout_17_rsc_rls_obj_iswt0),
      .dout_17_rsc_rls_obj_ld_core_sct(dout_17_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1 (
  clk, rst, tmp_17_data_rsci_addra_d, tmp_17_data_rsci_addrb_d, tmp_17_data_rsci_douta_d,
      tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_17_data_rsci_oswt, tmp_17_data_rsci_addra_d_core,
      tmp_17_data_rsci_addrb_d_core, tmp_17_data_rsci_douta_d_mxwt, tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_17_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_17_data_rsci_addra_d;
  output [7:0] tmp_17_data_rsci_addrb_d;
  input [63:0] tmp_17_data_rsci_douta_d;
  output tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_17_data_rsci_oswt;
  input [7:0] tmp_17_data_rsci_addra_d_core;
  input [7:0] tmp_17_data_rsci_addrb_d_core;
  output [15:0] tmp_17_data_rsci_douta_d_mxwt;
  input tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_17_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_17_data_rsci_biwt;
  wire tmp_17_data_rsci_bdwt;
  wire tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_17_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_17_data_rsci_addra_d_reg;
  wire tmp_17_data_rsci_biwt_iff;
  wire [7:0] tmp_17_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_dp_inst_tmp_17_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_dp_inst_tmp_17_data_rsci_addra_d_core
      = {1'b0 , (tmp_17_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_dp_inst_tmp_17_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_dp_inst_tmp_17_data_rsci_addrb_d_core
      = {1'b0 , (tmp_17_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_17_data_rsci_oswt(tmp_17_data_rsci_oswt),
      .tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_17_data_rsci_biwt(tmp_17_data_rsci_biwt),
      .tmp_17_data_rsci_bdwt(tmp_17_data_rsci_bdwt),
      .tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_17_data_rsci_biwt_pff(tmp_17_data_rsci_biwt_iff),
      .tmp_17_data_rsci_oswt_pff(tmp_17_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_17_data_rsci_addra_d(tmp_17_data_rsci_addra_d_reg),
      .tmp_17_data_rsci_addrb_d(tmp_17_data_rsci_addrb_d_reg),
      .tmp_17_data_rsci_douta_d(tmp_17_data_rsci_douta_d),
      .tmp_17_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_dp_inst_tmp_17_data_rsci_addra_d_core[7:0]),
      .tmp_17_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_tmp_17_data_rsc_wait_dp_inst_tmp_17_data_rsci_addrb_d_core[7:0]),
      .tmp_17_data_rsci_douta_d_mxwt(tmp_17_data_rsci_douta_d_mxwt_pconst),
      .tmp_17_data_rsci_biwt(tmp_17_data_rsci_biwt),
      .tmp_17_data_rsci_bdwt(tmp_17_data_rsci_bdwt),
      .tmp_17_data_rsci_biwt_pff(tmp_17_data_rsci_biwt_iff)
    );
  assign tmp_17_data_rsci_douta_d_mxwt = tmp_17_data_rsci_douta_d_mxwt_pconst;
  assign tmp_17_data_rsci_addra_d = tmp_17_data_rsci_addra_d_reg;
  assign tmp_17_data_rsci_addrb_d = tmp_17_data_rsci_addrb_d_reg;
  assign tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1 (
  clk, rst, tmp_16_data_rsci_addra_d, tmp_16_data_rsci_addrb_d, tmp_16_data_rsci_douta_d,
      tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_16_data_rsci_oswt, tmp_16_data_rsci_addra_d_core,
      tmp_16_data_rsci_addrb_d_core, tmp_16_data_rsci_douta_d_mxwt, tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_16_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_16_data_rsci_addra_d;
  output [7:0] tmp_16_data_rsci_addrb_d;
  input [63:0] tmp_16_data_rsci_douta_d;
  output tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_16_data_rsci_oswt;
  input [7:0] tmp_16_data_rsci_addra_d_core;
  input [7:0] tmp_16_data_rsci_addrb_d_core;
  output [15:0] tmp_16_data_rsci_douta_d_mxwt;
  input tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_16_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_16_data_rsci_biwt;
  wire tmp_16_data_rsci_bdwt;
  wire tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_16_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_16_data_rsci_addra_d_reg;
  wire tmp_16_data_rsci_biwt_iff;
  wire [7:0] tmp_16_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_dp_inst_tmp_16_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_dp_inst_tmp_16_data_rsci_addra_d_core
      = {1'b0 , (tmp_16_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_dp_inst_tmp_16_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_dp_inst_tmp_16_data_rsci_addrb_d_core
      = {1'b0 , (tmp_16_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_16_data_rsci_oswt(tmp_16_data_rsci_oswt),
      .tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_16_data_rsci_biwt(tmp_16_data_rsci_biwt),
      .tmp_16_data_rsci_bdwt(tmp_16_data_rsci_bdwt),
      .tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_16_data_rsci_biwt_pff(tmp_16_data_rsci_biwt_iff),
      .tmp_16_data_rsci_oswt_pff(tmp_16_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_16_data_rsci_addra_d(tmp_16_data_rsci_addra_d_reg),
      .tmp_16_data_rsci_addrb_d(tmp_16_data_rsci_addrb_d_reg),
      .tmp_16_data_rsci_douta_d(tmp_16_data_rsci_douta_d),
      .tmp_16_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_dp_inst_tmp_16_data_rsci_addra_d_core[7:0]),
      .tmp_16_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_tmp_16_data_rsc_wait_dp_inst_tmp_16_data_rsci_addrb_d_core[7:0]),
      .tmp_16_data_rsci_douta_d_mxwt(tmp_16_data_rsci_douta_d_mxwt_pconst),
      .tmp_16_data_rsci_biwt(tmp_16_data_rsci_biwt),
      .tmp_16_data_rsci_bdwt(tmp_16_data_rsci_bdwt),
      .tmp_16_data_rsci_biwt_pff(tmp_16_data_rsci_biwt_iff)
    );
  assign tmp_16_data_rsci_douta_d_mxwt = tmp_16_data_rsci_douta_d_mxwt_pconst;
  assign tmp_16_data_rsci_addra_d = tmp_16_data_rsci_addra_d_reg;
  assign tmp_16_data_rsci_addrb_d = tmp_16_data_rsci_addrb_d_reg;
  assign tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1 (
  clk, rst, tmp_15_data_rsci_addra_d, tmp_15_data_rsci_addrb_d, tmp_15_data_rsci_douta_d,
      tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_15_data_rsci_oswt, tmp_15_data_rsci_addra_d_core,
      tmp_15_data_rsci_addrb_d_core, tmp_15_data_rsci_douta_d_mxwt, tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_15_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_15_data_rsci_addra_d;
  output [7:0] tmp_15_data_rsci_addrb_d;
  input [63:0] tmp_15_data_rsci_douta_d;
  output tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_15_data_rsci_oswt;
  input [7:0] tmp_15_data_rsci_addra_d_core;
  input [7:0] tmp_15_data_rsci_addrb_d_core;
  output [15:0] tmp_15_data_rsci_douta_d_mxwt;
  input tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_15_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_15_data_rsci_biwt;
  wire tmp_15_data_rsci_bdwt;
  wire tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_15_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_15_data_rsci_addra_d_reg;
  wire tmp_15_data_rsci_biwt_iff;
  wire [7:0] tmp_15_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_dp_inst_tmp_15_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_dp_inst_tmp_15_data_rsci_addra_d_core
      = {1'b0 , (tmp_15_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_dp_inst_tmp_15_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_dp_inst_tmp_15_data_rsci_addrb_d_core
      = {1'b0 , (tmp_15_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_15_data_rsci_oswt(tmp_15_data_rsci_oswt),
      .tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_15_data_rsci_biwt(tmp_15_data_rsci_biwt),
      .tmp_15_data_rsci_bdwt(tmp_15_data_rsci_bdwt),
      .tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_15_data_rsci_biwt_pff(tmp_15_data_rsci_biwt_iff),
      .tmp_15_data_rsci_oswt_pff(tmp_15_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_15_data_rsci_addra_d(tmp_15_data_rsci_addra_d_reg),
      .tmp_15_data_rsci_addrb_d(tmp_15_data_rsci_addrb_d_reg),
      .tmp_15_data_rsci_douta_d(tmp_15_data_rsci_douta_d),
      .tmp_15_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_dp_inst_tmp_15_data_rsci_addra_d_core[7:0]),
      .tmp_15_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_tmp_15_data_rsc_wait_dp_inst_tmp_15_data_rsci_addrb_d_core[7:0]),
      .tmp_15_data_rsci_douta_d_mxwt(tmp_15_data_rsci_douta_d_mxwt_pconst),
      .tmp_15_data_rsci_biwt(tmp_15_data_rsci_biwt),
      .tmp_15_data_rsci_bdwt(tmp_15_data_rsci_bdwt),
      .tmp_15_data_rsci_biwt_pff(tmp_15_data_rsci_biwt_iff)
    );
  assign tmp_15_data_rsci_douta_d_mxwt = tmp_15_data_rsci_douta_d_mxwt_pconst;
  assign tmp_15_data_rsci_addra_d = tmp_15_data_rsci_addra_d_reg;
  assign tmp_15_data_rsci_addrb_d = tmp_15_data_rsci_addrb_d_reg;
  assign tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1 (
  clk, rst, tmp_14_data_rsci_addra_d, tmp_14_data_rsci_addrb_d, tmp_14_data_rsci_douta_d,
      tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_14_data_rsci_oswt, tmp_14_data_rsci_addra_d_core,
      tmp_14_data_rsci_addrb_d_core, tmp_14_data_rsci_douta_d_mxwt, tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_14_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_14_data_rsci_addra_d;
  output [7:0] tmp_14_data_rsci_addrb_d;
  input [63:0] tmp_14_data_rsci_douta_d;
  output tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_14_data_rsci_oswt;
  input [7:0] tmp_14_data_rsci_addra_d_core;
  input [7:0] tmp_14_data_rsci_addrb_d_core;
  output [15:0] tmp_14_data_rsci_douta_d_mxwt;
  input tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_14_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_14_data_rsci_biwt;
  wire tmp_14_data_rsci_bdwt;
  wire tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_14_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_14_data_rsci_addra_d_reg;
  wire tmp_14_data_rsci_biwt_iff;
  wire [7:0] tmp_14_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_dp_inst_tmp_14_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_dp_inst_tmp_14_data_rsci_addra_d_core
      = {1'b0 , (tmp_14_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_dp_inst_tmp_14_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_dp_inst_tmp_14_data_rsci_addrb_d_core
      = {1'b0 , (tmp_14_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_14_data_rsci_oswt(tmp_14_data_rsci_oswt),
      .tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_14_data_rsci_biwt(tmp_14_data_rsci_biwt),
      .tmp_14_data_rsci_bdwt(tmp_14_data_rsci_bdwt),
      .tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_14_data_rsci_biwt_pff(tmp_14_data_rsci_biwt_iff),
      .tmp_14_data_rsci_oswt_pff(tmp_14_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_14_data_rsci_addra_d(tmp_14_data_rsci_addra_d_reg),
      .tmp_14_data_rsci_addrb_d(tmp_14_data_rsci_addrb_d_reg),
      .tmp_14_data_rsci_douta_d(tmp_14_data_rsci_douta_d),
      .tmp_14_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_dp_inst_tmp_14_data_rsci_addra_d_core[7:0]),
      .tmp_14_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_tmp_14_data_rsc_wait_dp_inst_tmp_14_data_rsci_addrb_d_core[7:0]),
      .tmp_14_data_rsci_douta_d_mxwt(tmp_14_data_rsci_douta_d_mxwt_pconst),
      .tmp_14_data_rsci_biwt(tmp_14_data_rsci_biwt),
      .tmp_14_data_rsci_bdwt(tmp_14_data_rsci_bdwt),
      .tmp_14_data_rsci_biwt_pff(tmp_14_data_rsci_biwt_iff)
    );
  assign tmp_14_data_rsci_douta_d_mxwt = tmp_14_data_rsci_douta_d_mxwt_pconst;
  assign tmp_14_data_rsci_addra_d = tmp_14_data_rsci_addra_d_reg;
  assign tmp_14_data_rsci_addrb_d = tmp_14_data_rsci_addrb_d_reg;
  assign tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1 (
  clk, rst, tmp_13_data_rsci_addra_d, tmp_13_data_rsci_addrb_d, tmp_13_data_rsci_douta_d,
      tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_13_data_rsci_oswt, tmp_13_data_rsci_addra_d_core,
      tmp_13_data_rsci_addrb_d_core, tmp_13_data_rsci_douta_d_mxwt, tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_13_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_13_data_rsci_addra_d;
  output [7:0] tmp_13_data_rsci_addrb_d;
  input [63:0] tmp_13_data_rsci_douta_d;
  output tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_13_data_rsci_oswt;
  input [7:0] tmp_13_data_rsci_addra_d_core;
  input [7:0] tmp_13_data_rsci_addrb_d_core;
  output [15:0] tmp_13_data_rsci_douta_d_mxwt;
  input tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_13_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_13_data_rsci_biwt;
  wire tmp_13_data_rsci_bdwt;
  wire tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_13_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_13_data_rsci_addra_d_reg;
  wire tmp_13_data_rsci_biwt_iff;
  wire [7:0] tmp_13_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_dp_inst_tmp_13_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_dp_inst_tmp_13_data_rsci_addra_d_core
      = {1'b0 , (tmp_13_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_dp_inst_tmp_13_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_dp_inst_tmp_13_data_rsci_addrb_d_core
      = {1'b0 , (tmp_13_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_13_data_rsci_oswt(tmp_13_data_rsci_oswt),
      .tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_13_data_rsci_biwt(tmp_13_data_rsci_biwt),
      .tmp_13_data_rsci_bdwt(tmp_13_data_rsci_bdwt),
      .tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_13_data_rsci_biwt_pff(tmp_13_data_rsci_biwt_iff),
      .tmp_13_data_rsci_oswt_pff(tmp_13_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_13_data_rsci_addra_d(tmp_13_data_rsci_addra_d_reg),
      .tmp_13_data_rsci_addrb_d(tmp_13_data_rsci_addrb_d_reg),
      .tmp_13_data_rsci_douta_d(tmp_13_data_rsci_douta_d),
      .tmp_13_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_dp_inst_tmp_13_data_rsci_addra_d_core[7:0]),
      .tmp_13_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_tmp_13_data_rsc_wait_dp_inst_tmp_13_data_rsci_addrb_d_core[7:0]),
      .tmp_13_data_rsci_douta_d_mxwt(tmp_13_data_rsci_douta_d_mxwt_pconst),
      .tmp_13_data_rsci_biwt(tmp_13_data_rsci_biwt),
      .tmp_13_data_rsci_bdwt(tmp_13_data_rsci_bdwt),
      .tmp_13_data_rsci_biwt_pff(tmp_13_data_rsci_biwt_iff)
    );
  assign tmp_13_data_rsci_douta_d_mxwt = tmp_13_data_rsci_douta_d_mxwt_pconst;
  assign tmp_13_data_rsci_addra_d = tmp_13_data_rsci_addra_d_reg;
  assign tmp_13_data_rsci_addrb_d = tmp_13_data_rsci_addrb_d_reg;
  assign tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1 (
  clk, rst, tmp_12_data_rsci_addra_d, tmp_12_data_rsci_addrb_d, tmp_12_data_rsci_douta_d,
      tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_12_data_rsci_oswt, tmp_12_data_rsci_addra_d_core,
      tmp_12_data_rsci_addrb_d_core, tmp_12_data_rsci_douta_d_mxwt, tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_12_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_12_data_rsci_addra_d;
  output [7:0] tmp_12_data_rsci_addrb_d;
  input [63:0] tmp_12_data_rsci_douta_d;
  output tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_12_data_rsci_oswt;
  input [7:0] tmp_12_data_rsci_addra_d_core;
  input [7:0] tmp_12_data_rsci_addrb_d_core;
  output [15:0] tmp_12_data_rsci_douta_d_mxwt;
  input tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_12_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_12_data_rsci_biwt;
  wire tmp_12_data_rsci_bdwt;
  wire tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_12_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_12_data_rsci_addra_d_reg;
  wire tmp_12_data_rsci_biwt_iff;
  wire [7:0] tmp_12_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_dp_inst_tmp_12_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_dp_inst_tmp_12_data_rsci_addra_d_core
      = {1'b0 , (tmp_12_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_dp_inst_tmp_12_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_dp_inst_tmp_12_data_rsci_addrb_d_core
      = {1'b0 , (tmp_12_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_12_data_rsci_oswt(tmp_12_data_rsci_oswt),
      .tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_12_data_rsci_biwt(tmp_12_data_rsci_biwt),
      .tmp_12_data_rsci_bdwt(tmp_12_data_rsci_bdwt),
      .tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_12_data_rsci_biwt_pff(tmp_12_data_rsci_biwt_iff),
      .tmp_12_data_rsci_oswt_pff(tmp_12_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_12_data_rsci_addra_d(tmp_12_data_rsci_addra_d_reg),
      .tmp_12_data_rsci_addrb_d(tmp_12_data_rsci_addrb_d_reg),
      .tmp_12_data_rsci_douta_d(tmp_12_data_rsci_douta_d),
      .tmp_12_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_dp_inst_tmp_12_data_rsci_addra_d_core[7:0]),
      .tmp_12_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_tmp_12_data_rsc_wait_dp_inst_tmp_12_data_rsci_addrb_d_core[7:0]),
      .tmp_12_data_rsci_douta_d_mxwt(tmp_12_data_rsci_douta_d_mxwt_pconst),
      .tmp_12_data_rsci_biwt(tmp_12_data_rsci_biwt),
      .tmp_12_data_rsci_bdwt(tmp_12_data_rsci_bdwt),
      .tmp_12_data_rsci_biwt_pff(tmp_12_data_rsci_biwt_iff)
    );
  assign tmp_12_data_rsci_douta_d_mxwt = tmp_12_data_rsci_douta_d_mxwt_pconst;
  assign tmp_12_data_rsci_addra_d = tmp_12_data_rsci_addra_d_reg;
  assign tmp_12_data_rsci_addrb_d = tmp_12_data_rsci_addrb_d_reg;
  assign tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1 (
  clk, rst, tmp_11_data_rsci_addra_d, tmp_11_data_rsci_addrb_d, tmp_11_data_rsci_douta_d,
      tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_11_data_rsci_oswt, tmp_11_data_rsci_addra_d_core,
      tmp_11_data_rsci_addrb_d_core, tmp_11_data_rsci_douta_d_mxwt, tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_11_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_11_data_rsci_addra_d;
  output [7:0] tmp_11_data_rsci_addrb_d;
  input [63:0] tmp_11_data_rsci_douta_d;
  output tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_11_data_rsci_oswt;
  input [7:0] tmp_11_data_rsci_addra_d_core;
  input [7:0] tmp_11_data_rsci_addrb_d_core;
  output [15:0] tmp_11_data_rsci_douta_d_mxwt;
  input tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_11_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_11_data_rsci_biwt;
  wire tmp_11_data_rsci_bdwt;
  wire tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_11_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_11_data_rsci_addra_d_reg;
  wire tmp_11_data_rsci_biwt_iff;
  wire [7:0] tmp_11_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_dp_inst_tmp_11_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_dp_inst_tmp_11_data_rsci_addra_d_core
      = {1'b0 , (tmp_11_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_dp_inst_tmp_11_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_dp_inst_tmp_11_data_rsci_addrb_d_core
      = {1'b0 , (tmp_11_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_11_data_rsci_oswt(tmp_11_data_rsci_oswt),
      .tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_11_data_rsci_biwt(tmp_11_data_rsci_biwt),
      .tmp_11_data_rsci_bdwt(tmp_11_data_rsci_bdwt),
      .tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_11_data_rsci_biwt_pff(tmp_11_data_rsci_biwt_iff),
      .tmp_11_data_rsci_oswt_pff(tmp_11_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_11_data_rsci_addra_d(tmp_11_data_rsci_addra_d_reg),
      .tmp_11_data_rsci_addrb_d(tmp_11_data_rsci_addrb_d_reg),
      .tmp_11_data_rsci_douta_d(tmp_11_data_rsci_douta_d),
      .tmp_11_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_dp_inst_tmp_11_data_rsci_addra_d_core[7:0]),
      .tmp_11_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_tmp_11_data_rsc_wait_dp_inst_tmp_11_data_rsci_addrb_d_core[7:0]),
      .tmp_11_data_rsci_douta_d_mxwt(tmp_11_data_rsci_douta_d_mxwt_pconst),
      .tmp_11_data_rsci_biwt(tmp_11_data_rsci_biwt),
      .tmp_11_data_rsci_bdwt(tmp_11_data_rsci_bdwt),
      .tmp_11_data_rsci_biwt_pff(tmp_11_data_rsci_biwt_iff)
    );
  assign tmp_11_data_rsci_douta_d_mxwt = tmp_11_data_rsci_douta_d_mxwt_pconst;
  assign tmp_11_data_rsci_addra_d = tmp_11_data_rsci_addra_d_reg;
  assign tmp_11_data_rsci_addrb_d = tmp_11_data_rsci_addrb_d_reg;
  assign tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1 (
  clk, rst, tmp_10_data_rsci_addra_d, tmp_10_data_rsci_addrb_d, tmp_10_data_rsci_douta_d,
      tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_10_data_rsci_oswt, tmp_10_data_rsci_addra_d_core,
      tmp_10_data_rsci_addrb_d_core, tmp_10_data_rsci_douta_d_mxwt, tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_10_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_10_data_rsci_addra_d;
  output [7:0] tmp_10_data_rsci_addrb_d;
  input [63:0] tmp_10_data_rsci_douta_d;
  output tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_10_data_rsci_oswt;
  input [7:0] tmp_10_data_rsci_addra_d_core;
  input [7:0] tmp_10_data_rsci_addrb_d_core;
  output [15:0] tmp_10_data_rsci_douta_d_mxwt;
  input tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_10_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_10_data_rsci_biwt;
  wire tmp_10_data_rsci_bdwt;
  wire tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_10_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_10_data_rsci_addra_d_reg;
  wire tmp_10_data_rsci_biwt_iff;
  wire [7:0] tmp_10_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_dp_inst_tmp_10_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_dp_inst_tmp_10_data_rsci_addra_d_core
      = {1'b0 , (tmp_10_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_dp_inst_tmp_10_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_dp_inst_tmp_10_data_rsci_addrb_d_core
      = {1'b0 , (tmp_10_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_10_data_rsci_oswt(tmp_10_data_rsci_oswt),
      .tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_10_data_rsci_biwt(tmp_10_data_rsci_biwt),
      .tmp_10_data_rsci_bdwt(tmp_10_data_rsci_bdwt),
      .tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_10_data_rsci_biwt_pff(tmp_10_data_rsci_biwt_iff),
      .tmp_10_data_rsci_oswt_pff(tmp_10_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_10_data_rsci_addra_d(tmp_10_data_rsci_addra_d_reg),
      .tmp_10_data_rsci_addrb_d(tmp_10_data_rsci_addrb_d_reg),
      .tmp_10_data_rsci_douta_d(tmp_10_data_rsci_douta_d),
      .tmp_10_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_dp_inst_tmp_10_data_rsci_addra_d_core[7:0]),
      .tmp_10_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_tmp_10_data_rsc_wait_dp_inst_tmp_10_data_rsci_addrb_d_core[7:0]),
      .tmp_10_data_rsci_douta_d_mxwt(tmp_10_data_rsci_douta_d_mxwt_pconst),
      .tmp_10_data_rsci_biwt(tmp_10_data_rsci_biwt),
      .tmp_10_data_rsci_bdwt(tmp_10_data_rsci_bdwt),
      .tmp_10_data_rsci_biwt_pff(tmp_10_data_rsci_biwt_iff)
    );
  assign tmp_10_data_rsci_douta_d_mxwt = tmp_10_data_rsci_douta_d_mxwt_pconst;
  assign tmp_10_data_rsci_addra_d = tmp_10_data_rsci_addra_d_reg;
  assign tmp_10_data_rsci_addrb_d = tmp_10_data_rsci_addrb_d_reg;
  assign tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1 (
  clk, rst, tmp_9_data_rsci_addra_d, tmp_9_data_rsci_addrb_d, tmp_9_data_rsci_douta_d,
      tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_9_data_rsci_oswt, tmp_9_data_rsci_addra_d_core, tmp_9_data_rsci_addrb_d_core,
      tmp_9_data_rsci_douta_d_mxwt, tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_9_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_9_data_rsci_addra_d;
  output [7:0] tmp_9_data_rsci_addrb_d;
  input [63:0] tmp_9_data_rsci_douta_d;
  output tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_9_data_rsci_oswt;
  input [7:0] tmp_9_data_rsci_addra_d_core;
  input [7:0] tmp_9_data_rsci_addrb_d_core;
  output [15:0] tmp_9_data_rsci_douta_d_mxwt;
  input tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_9_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_9_data_rsci_biwt;
  wire tmp_9_data_rsci_bdwt;
  wire tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_9_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_9_data_rsci_addra_d_reg;
  wire tmp_9_data_rsci_biwt_iff;
  wire [7:0] tmp_9_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_dp_inst_tmp_9_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_dp_inst_tmp_9_data_rsci_addra_d_core
      = {1'b0 , (tmp_9_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_dp_inst_tmp_9_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_dp_inst_tmp_9_data_rsci_addrb_d_core
      = {1'b0 , (tmp_9_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_9_data_rsci_oswt(tmp_9_data_rsci_oswt),
      .tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_9_data_rsci_biwt(tmp_9_data_rsci_biwt),
      .tmp_9_data_rsci_bdwt(tmp_9_data_rsci_bdwt),
      .tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_9_data_rsci_biwt_pff(tmp_9_data_rsci_biwt_iff),
      .tmp_9_data_rsci_oswt_pff(tmp_9_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_9_data_rsci_addra_d(tmp_9_data_rsci_addra_d_reg),
      .tmp_9_data_rsci_addrb_d(tmp_9_data_rsci_addrb_d_reg),
      .tmp_9_data_rsci_douta_d(tmp_9_data_rsci_douta_d),
      .tmp_9_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_dp_inst_tmp_9_data_rsci_addra_d_core[7:0]),
      .tmp_9_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_tmp_9_data_rsc_wait_dp_inst_tmp_9_data_rsci_addrb_d_core[7:0]),
      .tmp_9_data_rsci_douta_d_mxwt(tmp_9_data_rsci_douta_d_mxwt_pconst),
      .tmp_9_data_rsci_biwt(tmp_9_data_rsci_biwt),
      .tmp_9_data_rsci_bdwt(tmp_9_data_rsci_bdwt),
      .tmp_9_data_rsci_biwt_pff(tmp_9_data_rsci_biwt_iff)
    );
  assign tmp_9_data_rsci_douta_d_mxwt = tmp_9_data_rsci_douta_d_mxwt_pconst;
  assign tmp_9_data_rsci_addra_d = tmp_9_data_rsci_addra_d_reg;
  assign tmp_9_data_rsci_addrb_d = tmp_9_data_rsci_addrb_d_reg;
  assign tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1 (
  clk, rst, tmp_8_data_rsci_addra_d, tmp_8_data_rsci_addrb_d, tmp_8_data_rsci_douta_d,
      tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_8_data_rsci_oswt, tmp_8_data_rsci_addra_d_core, tmp_8_data_rsci_addrb_d_core,
      tmp_8_data_rsci_douta_d_mxwt, tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_8_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_8_data_rsci_addra_d;
  output [7:0] tmp_8_data_rsci_addrb_d;
  input [63:0] tmp_8_data_rsci_douta_d;
  output tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_8_data_rsci_oswt;
  input [7:0] tmp_8_data_rsci_addra_d_core;
  input [7:0] tmp_8_data_rsci_addrb_d_core;
  output [15:0] tmp_8_data_rsci_douta_d_mxwt;
  input tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_8_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_8_data_rsci_biwt;
  wire tmp_8_data_rsci_bdwt;
  wire tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_8_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_8_data_rsci_addra_d_reg;
  wire tmp_8_data_rsci_biwt_iff;
  wire [7:0] tmp_8_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_dp_inst_tmp_8_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_dp_inst_tmp_8_data_rsci_addra_d_core
      = {1'b0 , (tmp_8_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_dp_inst_tmp_8_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_dp_inst_tmp_8_data_rsci_addrb_d_core
      = {1'b0 , (tmp_8_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_8_data_rsci_oswt(tmp_8_data_rsci_oswt),
      .tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_8_data_rsci_biwt(tmp_8_data_rsci_biwt),
      .tmp_8_data_rsci_bdwt(tmp_8_data_rsci_bdwt),
      .tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_8_data_rsci_biwt_pff(tmp_8_data_rsci_biwt_iff),
      .tmp_8_data_rsci_oswt_pff(tmp_8_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_8_data_rsci_addra_d(tmp_8_data_rsci_addra_d_reg),
      .tmp_8_data_rsci_addrb_d(tmp_8_data_rsci_addrb_d_reg),
      .tmp_8_data_rsci_douta_d(tmp_8_data_rsci_douta_d),
      .tmp_8_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_dp_inst_tmp_8_data_rsci_addra_d_core[7:0]),
      .tmp_8_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_tmp_8_data_rsc_wait_dp_inst_tmp_8_data_rsci_addrb_d_core[7:0]),
      .tmp_8_data_rsci_douta_d_mxwt(tmp_8_data_rsci_douta_d_mxwt_pconst),
      .tmp_8_data_rsci_biwt(tmp_8_data_rsci_biwt),
      .tmp_8_data_rsci_bdwt(tmp_8_data_rsci_bdwt),
      .tmp_8_data_rsci_biwt_pff(tmp_8_data_rsci_biwt_iff)
    );
  assign tmp_8_data_rsci_douta_d_mxwt = tmp_8_data_rsci_douta_d_mxwt_pconst;
  assign tmp_8_data_rsci_addra_d = tmp_8_data_rsci_addra_d_reg;
  assign tmp_8_data_rsci_addrb_d = tmp_8_data_rsci_addrb_d_reg;
  assign tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1 (
  clk, rst, tmp_7_data_rsci_addra_d, tmp_7_data_rsci_addrb_d, tmp_7_data_rsci_douta_d,
      tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_7_data_rsci_oswt, tmp_7_data_rsci_addra_d_core, tmp_7_data_rsci_addrb_d_core,
      tmp_7_data_rsci_douta_d_mxwt, tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_7_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_7_data_rsci_addra_d;
  output [7:0] tmp_7_data_rsci_addrb_d;
  input [63:0] tmp_7_data_rsci_douta_d;
  output tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_7_data_rsci_oswt;
  input [7:0] tmp_7_data_rsci_addra_d_core;
  input [7:0] tmp_7_data_rsci_addrb_d_core;
  output [15:0] tmp_7_data_rsci_douta_d_mxwt;
  input tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_7_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_7_data_rsci_biwt;
  wire tmp_7_data_rsci_bdwt;
  wire tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_7_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_7_data_rsci_addra_d_reg;
  wire tmp_7_data_rsci_biwt_iff;
  wire [7:0] tmp_7_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_dp_inst_tmp_7_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_dp_inst_tmp_7_data_rsci_addra_d_core
      = {1'b0 , (tmp_7_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_dp_inst_tmp_7_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_dp_inst_tmp_7_data_rsci_addrb_d_core
      = {1'b0 , (tmp_7_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_7_data_rsci_oswt(tmp_7_data_rsci_oswt),
      .tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_7_data_rsci_biwt(tmp_7_data_rsci_biwt),
      .tmp_7_data_rsci_bdwt(tmp_7_data_rsci_bdwt),
      .tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_7_data_rsci_biwt_pff(tmp_7_data_rsci_biwt_iff),
      .tmp_7_data_rsci_oswt_pff(tmp_7_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_7_data_rsci_addra_d(tmp_7_data_rsci_addra_d_reg),
      .tmp_7_data_rsci_addrb_d(tmp_7_data_rsci_addrb_d_reg),
      .tmp_7_data_rsci_douta_d(tmp_7_data_rsci_douta_d),
      .tmp_7_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_dp_inst_tmp_7_data_rsci_addra_d_core[7:0]),
      .tmp_7_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_tmp_7_data_rsc_wait_dp_inst_tmp_7_data_rsci_addrb_d_core[7:0]),
      .tmp_7_data_rsci_douta_d_mxwt(tmp_7_data_rsci_douta_d_mxwt_pconst),
      .tmp_7_data_rsci_biwt(tmp_7_data_rsci_biwt),
      .tmp_7_data_rsci_bdwt(tmp_7_data_rsci_bdwt),
      .tmp_7_data_rsci_biwt_pff(tmp_7_data_rsci_biwt_iff)
    );
  assign tmp_7_data_rsci_douta_d_mxwt = tmp_7_data_rsci_douta_d_mxwt_pconst;
  assign tmp_7_data_rsci_addra_d = tmp_7_data_rsci_addra_d_reg;
  assign tmp_7_data_rsci_addrb_d = tmp_7_data_rsci_addrb_d_reg;
  assign tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1 (
  clk, rst, tmp_6_data_rsci_addra_d, tmp_6_data_rsci_addrb_d, tmp_6_data_rsci_douta_d,
      tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_6_data_rsci_oswt, tmp_6_data_rsci_addra_d_core, tmp_6_data_rsci_addrb_d_core,
      tmp_6_data_rsci_douta_d_mxwt, tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_6_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_6_data_rsci_addra_d;
  output [7:0] tmp_6_data_rsci_addrb_d;
  input [63:0] tmp_6_data_rsci_douta_d;
  output tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_6_data_rsci_oswt;
  input [7:0] tmp_6_data_rsci_addra_d_core;
  input [7:0] tmp_6_data_rsci_addrb_d_core;
  output [15:0] tmp_6_data_rsci_douta_d_mxwt;
  input tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_6_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_6_data_rsci_biwt;
  wire tmp_6_data_rsci_bdwt;
  wire tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_6_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_6_data_rsci_addra_d_reg;
  wire tmp_6_data_rsci_biwt_iff;
  wire [7:0] tmp_6_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_dp_inst_tmp_6_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_dp_inst_tmp_6_data_rsci_addra_d_core
      = {1'b0 , (tmp_6_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_dp_inst_tmp_6_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_dp_inst_tmp_6_data_rsci_addrb_d_core
      = {1'b0 , (tmp_6_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_6_data_rsci_oswt(tmp_6_data_rsci_oswt),
      .tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_6_data_rsci_biwt(tmp_6_data_rsci_biwt),
      .tmp_6_data_rsci_bdwt(tmp_6_data_rsci_bdwt),
      .tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_6_data_rsci_biwt_pff(tmp_6_data_rsci_biwt_iff),
      .tmp_6_data_rsci_oswt_pff(tmp_6_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_6_data_rsci_addra_d(tmp_6_data_rsci_addra_d_reg),
      .tmp_6_data_rsci_addrb_d(tmp_6_data_rsci_addrb_d_reg),
      .tmp_6_data_rsci_douta_d(tmp_6_data_rsci_douta_d),
      .tmp_6_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_dp_inst_tmp_6_data_rsci_addra_d_core[7:0]),
      .tmp_6_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_tmp_6_data_rsc_wait_dp_inst_tmp_6_data_rsci_addrb_d_core[7:0]),
      .tmp_6_data_rsci_douta_d_mxwt(tmp_6_data_rsci_douta_d_mxwt_pconst),
      .tmp_6_data_rsci_biwt(tmp_6_data_rsci_biwt),
      .tmp_6_data_rsci_bdwt(tmp_6_data_rsci_bdwt),
      .tmp_6_data_rsci_biwt_pff(tmp_6_data_rsci_biwt_iff)
    );
  assign tmp_6_data_rsci_douta_d_mxwt = tmp_6_data_rsci_douta_d_mxwt_pconst;
  assign tmp_6_data_rsci_addra_d = tmp_6_data_rsci_addra_d_reg;
  assign tmp_6_data_rsci_addrb_d = tmp_6_data_rsci_addrb_d_reg;
  assign tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1 (
  clk, rst, tmp_5_data_rsci_addra_d, tmp_5_data_rsci_addrb_d, tmp_5_data_rsci_douta_d,
      tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_5_data_rsci_oswt, tmp_5_data_rsci_addra_d_core, tmp_5_data_rsci_addrb_d_core,
      tmp_5_data_rsci_douta_d_mxwt, tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_5_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_5_data_rsci_addra_d;
  output [7:0] tmp_5_data_rsci_addrb_d;
  input [63:0] tmp_5_data_rsci_douta_d;
  output tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_5_data_rsci_oswt;
  input [7:0] tmp_5_data_rsci_addra_d_core;
  input [7:0] tmp_5_data_rsci_addrb_d_core;
  output [15:0] tmp_5_data_rsci_douta_d_mxwt;
  input tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_5_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_5_data_rsci_biwt;
  wire tmp_5_data_rsci_bdwt;
  wire tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_5_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_5_data_rsci_addra_d_reg;
  wire tmp_5_data_rsci_biwt_iff;
  wire [7:0] tmp_5_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_dp_inst_tmp_5_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_dp_inst_tmp_5_data_rsci_addra_d_core
      = {1'b0 , (tmp_5_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_dp_inst_tmp_5_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_dp_inst_tmp_5_data_rsci_addrb_d_core
      = {1'b0 , (tmp_5_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_5_data_rsci_oswt(tmp_5_data_rsci_oswt),
      .tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_5_data_rsci_biwt(tmp_5_data_rsci_biwt),
      .tmp_5_data_rsci_bdwt(tmp_5_data_rsci_bdwt),
      .tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_5_data_rsci_biwt_pff(tmp_5_data_rsci_biwt_iff),
      .tmp_5_data_rsci_oswt_pff(tmp_5_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_5_data_rsci_addra_d(tmp_5_data_rsci_addra_d_reg),
      .tmp_5_data_rsci_addrb_d(tmp_5_data_rsci_addrb_d_reg),
      .tmp_5_data_rsci_douta_d(tmp_5_data_rsci_douta_d),
      .tmp_5_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_dp_inst_tmp_5_data_rsci_addra_d_core[7:0]),
      .tmp_5_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_tmp_5_data_rsc_wait_dp_inst_tmp_5_data_rsci_addrb_d_core[7:0]),
      .tmp_5_data_rsci_douta_d_mxwt(tmp_5_data_rsci_douta_d_mxwt_pconst),
      .tmp_5_data_rsci_biwt(tmp_5_data_rsci_biwt),
      .tmp_5_data_rsci_bdwt(tmp_5_data_rsci_bdwt),
      .tmp_5_data_rsci_biwt_pff(tmp_5_data_rsci_biwt_iff)
    );
  assign tmp_5_data_rsci_douta_d_mxwt = tmp_5_data_rsci_douta_d_mxwt_pconst;
  assign tmp_5_data_rsci_addra_d = tmp_5_data_rsci_addra_d_reg;
  assign tmp_5_data_rsci_addrb_d = tmp_5_data_rsci_addrb_d_reg;
  assign tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1 (
  clk, rst, tmp_4_data_rsci_addra_d, tmp_4_data_rsci_addrb_d, tmp_4_data_rsci_douta_d,
      tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_4_data_rsci_oswt, tmp_4_data_rsci_addra_d_core, tmp_4_data_rsci_addrb_d_core,
      tmp_4_data_rsci_douta_d_mxwt, tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_4_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_4_data_rsci_addra_d;
  output [7:0] tmp_4_data_rsci_addrb_d;
  input [63:0] tmp_4_data_rsci_douta_d;
  output tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_4_data_rsci_oswt;
  input [7:0] tmp_4_data_rsci_addra_d_core;
  input [7:0] tmp_4_data_rsci_addrb_d_core;
  output [15:0] tmp_4_data_rsci_douta_d_mxwt;
  input tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_4_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_4_data_rsci_biwt;
  wire tmp_4_data_rsci_bdwt;
  wire tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_4_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_4_data_rsci_addra_d_reg;
  wire tmp_4_data_rsci_biwt_iff;
  wire [7:0] tmp_4_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_dp_inst_tmp_4_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_dp_inst_tmp_4_data_rsci_addra_d_core
      = {1'b0 , (tmp_4_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_dp_inst_tmp_4_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_dp_inst_tmp_4_data_rsci_addrb_d_core
      = {1'b0 , (tmp_4_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_4_data_rsci_oswt(tmp_4_data_rsci_oswt),
      .tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_4_data_rsci_biwt(tmp_4_data_rsci_biwt),
      .tmp_4_data_rsci_bdwt(tmp_4_data_rsci_bdwt),
      .tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_4_data_rsci_biwt_pff(tmp_4_data_rsci_biwt_iff),
      .tmp_4_data_rsci_oswt_pff(tmp_4_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_4_data_rsci_addra_d(tmp_4_data_rsci_addra_d_reg),
      .tmp_4_data_rsci_addrb_d(tmp_4_data_rsci_addrb_d_reg),
      .tmp_4_data_rsci_douta_d(tmp_4_data_rsci_douta_d),
      .tmp_4_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_dp_inst_tmp_4_data_rsci_addra_d_core[7:0]),
      .tmp_4_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_tmp_4_data_rsc_wait_dp_inst_tmp_4_data_rsci_addrb_d_core[7:0]),
      .tmp_4_data_rsci_douta_d_mxwt(tmp_4_data_rsci_douta_d_mxwt_pconst),
      .tmp_4_data_rsci_biwt(tmp_4_data_rsci_biwt),
      .tmp_4_data_rsci_bdwt(tmp_4_data_rsci_bdwt),
      .tmp_4_data_rsci_biwt_pff(tmp_4_data_rsci_biwt_iff)
    );
  assign tmp_4_data_rsci_douta_d_mxwt = tmp_4_data_rsci_douta_d_mxwt_pconst;
  assign tmp_4_data_rsci_addra_d = tmp_4_data_rsci_addra_d_reg;
  assign tmp_4_data_rsci_addrb_d = tmp_4_data_rsci_addrb_d_reg;
  assign tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1 (
  clk, rst, tmp_3_data_rsci_addra_d, tmp_3_data_rsci_addrb_d, tmp_3_data_rsci_douta_d,
      tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_3_data_rsci_oswt, tmp_3_data_rsci_addra_d_core, tmp_3_data_rsci_addrb_d_core,
      tmp_3_data_rsci_douta_d_mxwt, tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_3_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_3_data_rsci_addra_d;
  output [7:0] tmp_3_data_rsci_addrb_d;
  input [63:0] tmp_3_data_rsci_douta_d;
  output tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_3_data_rsci_oswt;
  input [7:0] tmp_3_data_rsci_addra_d_core;
  input [7:0] tmp_3_data_rsci_addrb_d_core;
  output [15:0] tmp_3_data_rsci_douta_d_mxwt;
  input tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_3_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_3_data_rsci_biwt;
  wire tmp_3_data_rsci_bdwt;
  wire tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_3_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_3_data_rsci_addra_d_reg;
  wire tmp_3_data_rsci_biwt_iff;
  wire [7:0] tmp_3_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_dp_inst_tmp_3_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_dp_inst_tmp_3_data_rsci_addra_d_core
      = {1'b0 , (tmp_3_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_dp_inst_tmp_3_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_dp_inst_tmp_3_data_rsci_addrb_d_core
      = {1'b0 , (tmp_3_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_3_data_rsci_oswt(tmp_3_data_rsci_oswt),
      .tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_3_data_rsci_biwt(tmp_3_data_rsci_biwt),
      .tmp_3_data_rsci_bdwt(tmp_3_data_rsci_bdwt),
      .tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_3_data_rsci_biwt_pff(tmp_3_data_rsci_biwt_iff),
      .tmp_3_data_rsci_oswt_pff(tmp_3_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_3_data_rsci_addra_d(tmp_3_data_rsci_addra_d_reg),
      .tmp_3_data_rsci_addrb_d(tmp_3_data_rsci_addrb_d_reg),
      .tmp_3_data_rsci_douta_d(tmp_3_data_rsci_douta_d),
      .tmp_3_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_dp_inst_tmp_3_data_rsci_addra_d_core[7:0]),
      .tmp_3_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_tmp_3_data_rsc_wait_dp_inst_tmp_3_data_rsci_addrb_d_core[7:0]),
      .tmp_3_data_rsci_douta_d_mxwt(tmp_3_data_rsci_douta_d_mxwt_pconst),
      .tmp_3_data_rsci_biwt(tmp_3_data_rsci_biwt),
      .tmp_3_data_rsci_bdwt(tmp_3_data_rsci_bdwt),
      .tmp_3_data_rsci_biwt_pff(tmp_3_data_rsci_biwt_iff)
    );
  assign tmp_3_data_rsci_douta_d_mxwt = tmp_3_data_rsci_douta_d_mxwt_pconst;
  assign tmp_3_data_rsci_addra_d = tmp_3_data_rsci_addra_d_reg;
  assign tmp_3_data_rsci_addrb_d = tmp_3_data_rsci_addrb_d_reg;
  assign tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1 (
  clk, rst, tmp_2_data_rsci_addra_d, tmp_2_data_rsci_addrb_d, tmp_2_data_rsci_douta_d,
      tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_2_data_rsci_oswt, tmp_2_data_rsci_addra_d_core, tmp_2_data_rsci_addrb_d_core,
      tmp_2_data_rsci_douta_d_mxwt, tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_2_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_2_data_rsci_addra_d;
  output [7:0] tmp_2_data_rsci_addrb_d;
  input [63:0] tmp_2_data_rsci_douta_d;
  output tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_2_data_rsci_oswt;
  input [7:0] tmp_2_data_rsci_addra_d_core;
  input [7:0] tmp_2_data_rsci_addrb_d_core;
  output [15:0] tmp_2_data_rsci_douta_d_mxwt;
  input tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_2_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_2_data_rsci_biwt;
  wire tmp_2_data_rsci_bdwt;
  wire tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_2_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_2_data_rsci_addra_d_reg;
  wire tmp_2_data_rsci_biwt_iff;
  wire [7:0] tmp_2_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_dp_inst_tmp_2_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_dp_inst_tmp_2_data_rsci_addra_d_core
      = {1'b0 , (tmp_2_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_dp_inst_tmp_2_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_dp_inst_tmp_2_data_rsci_addrb_d_core
      = {1'b0 , (tmp_2_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_2_data_rsci_oswt(tmp_2_data_rsci_oswt),
      .tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_2_data_rsci_biwt(tmp_2_data_rsci_biwt),
      .tmp_2_data_rsci_bdwt(tmp_2_data_rsci_bdwt),
      .tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_2_data_rsci_biwt_pff(tmp_2_data_rsci_biwt_iff),
      .tmp_2_data_rsci_oswt_pff(tmp_2_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_2_data_rsci_addra_d(tmp_2_data_rsci_addra_d_reg),
      .tmp_2_data_rsci_addrb_d(tmp_2_data_rsci_addrb_d_reg),
      .tmp_2_data_rsci_douta_d(tmp_2_data_rsci_douta_d),
      .tmp_2_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_dp_inst_tmp_2_data_rsci_addra_d_core[7:0]),
      .tmp_2_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_tmp_2_data_rsc_wait_dp_inst_tmp_2_data_rsci_addrb_d_core[7:0]),
      .tmp_2_data_rsci_douta_d_mxwt(tmp_2_data_rsci_douta_d_mxwt_pconst),
      .tmp_2_data_rsci_biwt(tmp_2_data_rsci_biwt),
      .tmp_2_data_rsci_bdwt(tmp_2_data_rsci_bdwt),
      .tmp_2_data_rsci_biwt_pff(tmp_2_data_rsci_biwt_iff)
    );
  assign tmp_2_data_rsci_douta_d_mxwt = tmp_2_data_rsci_douta_d_mxwt_pconst;
  assign tmp_2_data_rsci_addra_d = tmp_2_data_rsci_addra_d_reg;
  assign tmp_2_data_rsci_addrb_d = tmp_2_data_rsci_addrb_d_reg;
  assign tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1 (
  clk, rst, tmp_1_data_rsci_addra_d, tmp_1_data_rsci_addrb_d, tmp_1_data_rsci_douta_d,
      tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_1_data_rsci_oswt, tmp_1_data_rsci_addra_d_core, tmp_1_data_rsci_addrb_d_core,
      tmp_1_data_rsci_douta_d_mxwt, tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_1_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_1_data_rsci_addra_d;
  output [7:0] tmp_1_data_rsci_addrb_d;
  input [63:0] tmp_1_data_rsci_douta_d;
  output tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_1_data_rsci_oswt;
  input [7:0] tmp_1_data_rsci_addra_d_core;
  input [7:0] tmp_1_data_rsci_addrb_d_core;
  output [15:0] tmp_1_data_rsci_douta_d_mxwt;
  input tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_1_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_1_data_rsci_biwt;
  wire tmp_1_data_rsci_bdwt;
  wire tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_1_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_1_data_rsci_addra_d_reg;
  wire tmp_1_data_rsci_biwt_iff;
  wire [7:0] tmp_1_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_dp_inst_tmp_1_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_dp_inst_tmp_1_data_rsci_addra_d_core
      = {1'b0 , (tmp_1_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_dp_inst_tmp_1_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_dp_inst_tmp_1_data_rsci_addrb_d_core
      = {1'b0 , (tmp_1_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_1_data_rsci_oswt(tmp_1_data_rsci_oswt),
      .tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_1_data_rsci_biwt(tmp_1_data_rsci_biwt),
      .tmp_1_data_rsci_bdwt(tmp_1_data_rsci_bdwt),
      .tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_1_data_rsci_biwt_pff(tmp_1_data_rsci_biwt_iff),
      .tmp_1_data_rsci_oswt_pff(tmp_1_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_1_data_rsci_addra_d(tmp_1_data_rsci_addra_d_reg),
      .tmp_1_data_rsci_addrb_d(tmp_1_data_rsci_addrb_d_reg),
      .tmp_1_data_rsci_douta_d(tmp_1_data_rsci_douta_d),
      .tmp_1_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_dp_inst_tmp_1_data_rsci_addra_d_core[7:0]),
      .tmp_1_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_tmp_1_data_rsc_wait_dp_inst_tmp_1_data_rsci_addrb_d_core[7:0]),
      .tmp_1_data_rsci_douta_d_mxwt(tmp_1_data_rsci_douta_d_mxwt_pconst),
      .tmp_1_data_rsci_biwt(tmp_1_data_rsci_biwt),
      .tmp_1_data_rsci_bdwt(tmp_1_data_rsci_bdwt),
      .tmp_1_data_rsci_biwt_pff(tmp_1_data_rsci_biwt_iff)
    );
  assign tmp_1_data_rsci_douta_d_mxwt = tmp_1_data_rsci_douta_d_mxwt_pconst;
  assign tmp_1_data_rsci_addra_d = tmp_1_data_rsci_addra_d_reg;
  assign tmp_1_data_rsci_addrb_d = tmp_1_data_rsci_addrb_d_reg;
  assign tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1 (
  clk, rst, tmp_0_data_rsci_addra_d, tmp_0_data_rsci_addrb_d, tmp_0_data_rsci_douta_d,
      tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      core_wen, core_wten, tmp_0_data_rsci_oswt, tmp_0_data_rsci_addra_d_core, tmp_0_data_rsci_addrb_d_core,
      tmp_0_data_rsci_douta_d_mxwt, tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct,
      tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct, tmp_0_data_rsci_oswt_pff
);
  input clk;
  input rst;
  output [7:0] tmp_0_data_rsci_addra_d;
  output [7:0] tmp_0_data_rsci_addrb_d;
  input [63:0] tmp_0_data_rsci_douta_d;
  output tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wen;
  input core_wten;
  input tmp_0_data_rsci_oswt;
  input [7:0] tmp_0_data_rsci_addra_d_core;
  input [7:0] tmp_0_data_rsci_addrb_d_core;
  output [15:0] tmp_0_data_rsci_douta_d_mxwt;
  input tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  input tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  input tmp_0_data_rsci_oswt_pff;


  // Interconnect Declarations
  wire tmp_0_data_rsci_biwt;
  wire tmp_0_data_rsci_bdwt;
  wire tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  wire tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
  wire [15:0] tmp_0_data_rsci_douta_d_mxwt_pconst;
  wire [7:0] tmp_0_data_rsci_addra_d_reg;
  wire tmp_0_data_rsci_biwt_iff;
  wire [7:0] tmp_0_data_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_dp_inst_tmp_0_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_dp_inst_tmp_0_data_rsci_addra_d_core
      = {1'b0 , (tmp_0_data_rsci_addra_d_core[6:0])};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_dp_inst_tmp_0_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_dp_inst_tmp_0_data_rsci_addrb_d_core
      = {1'b0 , (tmp_0_data_rsci_addrb_d_core[6:0])};
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_ctrl
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_0_data_rsci_oswt(tmp_0_data_rsci_oswt),
      .tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct),
      .tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct),
      .tmp_0_data_rsci_biwt(tmp_0_data_rsci_biwt),
      .tmp_0_data_rsci_bdwt(tmp_0_data_rsci_bdwt),
      .tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct(tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct),
      .tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct),
      .tmp_0_data_rsci_biwt_pff(tmp_0_data_rsci_biwt_iff),
      .tmp_0_data_rsci_oswt_pff(tmp_0_data_rsci_oswt_pff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_dp
      WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_0_data_rsci_addra_d(tmp_0_data_rsci_addra_d_reg),
      .tmp_0_data_rsci_addrb_d(tmp_0_data_rsci_addrb_d_reg),
      .tmp_0_data_rsci_douta_d(tmp_0_data_rsci_douta_d),
      .tmp_0_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_dp_inst_tmp_0_data_rsci_addra_d_core[7:0]),
      .tmp_0_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_tmp_0_data_rsc_wait_dp_inst_tmp_0_data_rsci_addrb_d_core[7:0]),
      .tmp_0_data_rsci_douta_d_mxwt(tmp_0_data_rsci_douta_d_mxwt_pconst),
      .tmp_0_data_rsci_biwt(tmp_0_data_rsci_biwt),
      .tmp_0_data_rsci_bdwt(tmp_0_data_rsci_bdwt),
      .tmp_0_data_rsci_biwt_pff(tmp_0_data_rsci_biwt_iff)
    );
  assign tmp_0_data_rsci_douta_d_mxwt = tmp_0_data_rsci_douta_d_mxwt_pconst;
  assign tmp_0_data_rsci_addra_d = tmp_0_data_rsci_addra_d_reg;
  assign tmp_0_data_rsci_addrb_d = tmp_0_data_rsci_addrb_d_reg;
  assign tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_sct;
  assign tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1 (
  dout_17_rsci_dinb_d, dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_17_rsci_dinb_d_core,
      dout_17_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_17_rsci_dinb_d;
  output dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_17_rsci_dinb_d_core;
  input dout_17_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_17_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_dout_17_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_dout_17_rsc_wait_ctrl_inst
      (
      .dout_17_rsci_dinb_d_core_sct_pff(dout_17_rsci_dinb_d_core_sct_iff),
      .dout_17_rsci_iswt0_pff(dout_17_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_17_rsci_dinb_d = {(~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (~ dout_17_rsci_dinb_d_core_sct_iff) , (~ dout_17_rsci_dinb_d_core_sct_iff)
      , (dout_17_rsci_dinb_d_core[15:0])};
  assign dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_17_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1 (
  dout_16_rsci_dinb_d, dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_16_rsci_dinb_d_core,
      dout_16_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_16_rsci_dinb_d;
  output dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_16_rsci_dinb_d_core;
  input dout_16_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_16_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_dout_16_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_dout_16_rsc_wait_ctrl_inst
      (
      .dout_16_rsci_dinb_d_core_sct_pff(dout_16_rsci_dinb_d_core_sct_iff),
      .dout_16_rsci_iswt0_pff(dout_16_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_16_rsci_dinb_d = {(~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (~ dout_16_rsci_dinb_d_core_sct_iff) , (~ dout_16_rsci_dinb_d_core_sct_iff)
      , (dout_16_rsci_dinb_d_core[15:0])};
  assign dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_16_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1 (
  dout_15_rsci_dinb_d, dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_15_rsci_dinb_d_core,
      dout_15_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_15_rsci_dinb_d;
  output dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_15_rsci_dinb_d_core;
  input dout_15_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_15_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_dout_15_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_dout_15_rsc_wait_ctrl_inst
      (
      .dout_15_rsci_dinb_d_core_sct_pff(dout_15_rsci_dinb_d_core_sct_iff),
      .dout_15_rsci_iswt0_pff(dout_15_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_15_rsci_dinb_d = {(~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (~ dout_15_rsci_dinb_d_core_sct_iff) , (~ dout_15_rsci_dinb_d_core_sct_iff)
      , (dout_15_rsci_dinb_d_core[15:0])};
  assign dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_15_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1 (
  dout_14_rsci_dinb_d, dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_14_rsci_dinb_d_core,
      dout_14_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_14_rsci_dinb_d;
  output dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_14_rsci_dinb_d_core;
  input dout_14_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_14_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_dout_14_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_dout_14_rsc_wait_ctrl_inst
      (
      .dout_14_rsci_dinb_d_core_sct_pff(dout_14_rsci_dinb_d_core_sct_iff),
      .dout_14_rsci_iswt0_pff(dout_14_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_14_rsci_dinb_d = {(~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (~ dout_14_rsci_dinb_d_core_sct_iff) , (~ dout_14_rsci_dinb_d_core_sct_iff)
      , (dout_14_rsci_dinb_d_core[15:0])};
  assign dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_14_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1 (
  dout_13_rsci_dinb_d, dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_13_rsci_dinb_d_core,
      dout_13_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_13_rsci_dinb_d;
  output dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_13_rsci_dinb_d_core;
  input dout_13_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_13_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_dout_13_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_dout_13_rsc_wait_ctrl_inst
      (
      .dout_13_rsci_dinb_d_core_sct_pff(dout_13_rsci_dinb_d_core_sct_iff),
      .dout_13_rsci_iswt0_pff(dout_13_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_13_rsci_dinb_d = {(~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (~ dout_13_rsci_dinb_d_core_sct_iff) , (~ dout_13_rsci_dinb_d_core_sct_iff)
      , (dout_13_rsci_dinb_d_core[15:0])};
  assign dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_13_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1 (
  dout_12_rsci_dinb_d, dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_12_rsci_dinb_d_core,
      dout_12_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_12_rsci_dinb_d;
  output dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_12_rsci_dinb_d_core;
  input dout_12_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_12_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_dout_12_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_dout_12_rsc_wait_ctrl_inst
      (
      .dout_12_rsci_dinb_d_core_sct_pff(dout_12_rsci_dinb_d_core_sct_iff),
      .dout_12_rsci_iswt0_pff(dout_12_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_12_rsci_dinb_d = {(~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (~ dout_12_rsci_dinb_d_core_sct_iff) , (~ dout_12_rsci_dinb_d_core_sct_iff)
      , (dout_12_rsci_dinb_d_core[15:0])};
  assign dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_12_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1 (
  dout_11_rsci_dinb_d, dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_11_rsci_dinb_d_core,
      dout_11_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_11_rsci_dinb_d;
  output dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_11_rsci_dinb_d_core;
  input dout_11_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_11_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_dout_11_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_dout_11_rsc_wait_ctrl_inst
      (
      .dout_11_rsci_dinb_d_core_sct_pff(dout_11_rsci_dinb_d_core_sct_iff),
      .dout_11_rsci_iswt0_pff(dout_11_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_11_rsci_dinb_d = {(~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (~ dout_11_rsci_dinb_d_core_sct_iff) , (~ dout_11_rsci_dinb_d_core_sct_iff)
      , (dout_11_rsci_dinb_d_core[15:0])};
  assign dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_11_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1 (
  dout_10_rsci_dinb_d, dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_10_rsci_dinb_d_core,
      dout_10_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_10_rsci_dinb_d;
  output dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_10_rsci_dinb_d_core;
  input dout_10_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_10_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_dout_10_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_dout_10_rsc_wait_ctrl_inst
      (
      .dout_10_rsci_dinb_d_core_sct_pff(dout_10_rsci_dinb_d_core_sct_iff),
      .dout_10_rsci_iswt0_pff(dout_10_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_10_rsci_dinb_d = {(~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (~ dout_10_rsci_dinb_d_core_sct_iff) , (~ dout_10_rsci_dinb_d_core_sct_iff)
      , (dout_10_rsci_dinb_d_core[15:0])};
  assign dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_10_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1 (
  dout_9_rsci_dinb_d, dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_9_rsci_dinb_d_core,
      dout_9_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_9_rsci_dinb_d;
  output dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_9_rsci_dinb_d_core;
  input dout_9_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_9_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_dout_9_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_dout_9_rsc_wait_ctrl_inst
      (
      .dout_9_rsci_dinb_d_core_sct_pff(dout_9_rsci_dinb_d_core_sct_iff),
      .dout_9_rsci_iswt0_pff(dout_9_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_9_rsci_dinb_d = {(~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (~ dout_9_rsci_dinb_d_core_sct_iff) , (~ dout_9_rsci_dinb_d_core_sct_iff)
      , (dout_9_rsci_dinb_d_core[15:0])};
  assign dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_9_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1 (
  dout_8_rsci_dinb_d, dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_8_rsci_dinb_d_core,
      dout_8_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_8_rsci_dinb_d;
  output dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_8_rsci_dinb_d_core;
  input dout_8_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_8_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_dout_8_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_dout_8_rsc_wait_ctrl_inst
      (
      .dout_8_rsci_dinb_d_core_sct_pff(dout_8_rsci_dinb_d_core_sct_iff),
      .dout_8_rsci_iswt0_pff(dout_8_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_8_rsci_dinb_d = {(~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (~ dout_8_rsci_dinb_d_core_sct_iff) , (~ dout_8_rsci_dinb_d_core_sct_iff)
      , (dout_8_rsci_dinb_d_core[15:0])};
  assign dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_8_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1 (
  dout_7_rsci_dinb_d, dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_7_rsci_dinb_d_core,
      dout_7_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_7_rsci_dinb_d;
  output dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_7_rsci_dinb_d_core;
  input dout_7_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_7_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_dout_7_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_dout_7_rsc_wait_ctrl_inst
      (
      .dout_7_rsci_dinb_d_core_sct_pff(dout_7_rsci_dinb_d_core_sct_iff),
      .dout_7_rsci_iswt0_pff(dout_7_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_7_rsci_dinb_d = {(~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (~ dout_7_rsci_dinb_d_core_sct_iff) , (~ dout_7_rsci_dinb_d_core_sct_iff)
      , (dout_7_rsci_dinb_d_core[15:0])};
  assign dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_7_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1 (
  dout_6_rsci_dinb_d, dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_6_rsci_dinb_d_core,
      dout_6_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_6_rsci_dinb_d;
  output dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_6_rsci_dinb_d_core;
  input dout_6_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_6_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_dout_6_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_dout_6_rsc_wait_ctrl_inst
      (
      .dout_6_rsci_dinb_d_core_sct_pff(dout_6_rsci_dinb_d_core_sct_iff),
      .dout_6_rsci_iswt0_pff(dout_6_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_6_rsci_dinb_d = {(~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (~ dout_6_rsci_dinb_d_core_sct_iff) , (~ dout_6_rsci_dinb_d_core_sct_iff)
      , (dout_6_rsci_dinb_d_core[15:0])};
  assign dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_6_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1 (
  dout_5_rsci_dinb_d, dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_5_rsci_dinb_d_core,
      dout_5_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_5_rsci_dinb_d;
  output dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_5_rsci_dinb_d_core;
  input dout_5_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_5_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_dout_5_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_dout_5_rsc_wait_ctrl_inst
      (
      .dout_5_rsci_dinb_d_core_sct_pff(dout_5_rsci_dinb_d_core_sct_iff),
      .dout_5_rsci_iswt0_pff(dout_5_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_5_rsci_dinb_d = {(~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (~ dout_5_rsci_dinb_d_core_sct_iff) , (~ dout_5_rsci_dinb_d_core_sct_iff)
      , (dout_5_rsci_dinb_d_core[15:0])};
  assign dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_5_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1 (
  dout_4_rsci_dinb_d, dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_4_rsci_dinb_d_core,
      dout_4_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_4_rsci_dinb_d;
  output dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_4_rsci_dinb_d_core;
  input dout_4_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_4_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_dout_4_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_dout_4_rsc_wait_ctrl_inst
      (
      .dout_4_rsci_dinb_d_core_sct_pff(dout_4_rsci_dinb_d_core_sct_iff),
      .dout_4_rsci_iswt0_pff(dout_4_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_4_rsci_dinb_d = {(~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (~ dout_4_rsci_dinb_d_core_sct_iff) , (~ dout_4_rsci_dinb_d_core_sct_iff)
      , (dout_4_rsci_dinb_d_core[15:0])};
  assign dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_4_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1 (
  dout_3_rsci_dinb_d, dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_3_rsci_dinb_d_core,
      dout_3_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_3_rsci_dinb_d;
  output dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_3_rsci_dinb_d_core;
  input dout_3_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_3_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_dout_3_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_dout_3_rsc_wait_ctrl_inst
      (
      .dout_3_rsci_dinb_d_core_sct_pff(dout_3_rsci_dinb_d_core_sct_iff),
      .dout_3_rsci_iswt0_pff(dout_3_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_3_rsci_dinb_d = {(~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (~ dout_3_rsci_dinb_d_core_sct_iff) , (~ dout_3_rsci_dinb_d_core_sct_iff)
      , (dout_3_rsci_dinb_d_core[15:0])};
  assign dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_3_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1 (
  dout_2_rsci_dinb_d, dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_2_rsci_dinb_d_core,
      dout_2_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_2_rsci_dinb_d;
  output dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_2_rsci_dinb_d_core;
  input dout_2_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_2_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_dout_2_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_dout_2_rsc_wait_ctrl_inst
      (
      .dout_2_rsci_dinb_d_core_sct_pff(dout_2_rsci_dinb_d_core_sct_iff),
      .dout_2_rsci_iswt0_pff(dout_2_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_2_rsci_dinb_d = {(~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (~ dout_2_rsci_dinb_d_core_sct_iff) , (~ dout_2_rsci_dinb_d_core_sct_iff)
      , (dout_2_rsci_dinb_d_core[15:0])};
  assign dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_2_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1 (
  dout_1_rsci_dinb_d, dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_1_rsci_dinb_d_core,
      dout_1_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_1_rsci_dinb_d;
  output dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_1_rsci_dinb_d_core;
  input dout_1_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_1_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_dout_1_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_dout_1_rsc_wait_ctrl_inst
      (
      .dout_1_rsci_dinb_d_core_sct_pff(dout_1_rsci_dinb_d_core_sct_iff),
      .dout_1_rsci_iswt0_pff(dout_1_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_1_rsci_dinb_d = {(~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (~ dout_1_rsci_dinb_d_core_sct_iff) , (~ dout_1_rsci_dinb_d_core_sct_iff)
      , (dout_1_rsci_dinb_d_core[15:0])};
  assign dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_1_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1 (
  dout_0_rsci_dinb_d, dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_0_rsci_dinb_d_core,
      dout_0_rsci_iswt0_pff, core_wten_pff
);
  output [63:0] dout_0_rsci_dinb_d;
  output dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [63:0] dout_0_rsci_dinb_d_core;
  input dout_0_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_0_rsci_dinb_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_dout_0_rsc_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_dout_0_rsc_wait_ctrl_inst
      (
      .dout_0_rsci_dinb_d_core_sct_pff(dout_0_rsci_dinb_d_core_sct_iff),
      .dout_0_rsci_iswt0_pff(dout_0_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_0_rsci_dinb_d = {(~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (~ dout_0_rsci_dinb_d_core_sct_iff) , (~ dout_0_rsci_dinb_d_core_sct_iff)
      , (dout_0_rsci_dinb_d_core[15:0])};
  assign dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_0_rsci_dinb_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, core_wen, din_rsci_oswt, din_rsci_wen_comp,
      din_rsci_d_mxwt, core_wten
);
  input clk;
  input rst;
  input [15:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  input core_wen;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [15:0] din_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire din_rsci_ld_core_sct;
  wire din_rsci_vd;
  wire [15:0] din_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd16)) din_rsci (
      .ld(din_rsci_ld_core_sct),
      .vd(din_rsci_vd),
      .d(din_rsci_d),
      .lz(din_rsc_lz),
      .vz(din_rsc_vz),
      .z(din_rsc_z)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci_din_wait_ctrl WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci_din_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .din_rsci_oswt(din_rsci_oswt),
      .core_wten(core_wten),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_ld_core_sct(din_rsci_ld_core_sct),
      .din_rsci_vd(din_rsci_vd)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci_din_wait_dp WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci_din_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_d_mxwt(din_rsci_d_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_d(din_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj (
  clk, rst, din_0_rsc_req_vz, core_wen, core_wten, din_0_rsc_req_obj_oswt, din_0_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_0_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_0_rsc_req_obj_oswt;
  output din_0_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_0_rsc_req_obj_vd;
  wire din_0_rsc_req_obj_biwt;
  wire din_0_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_0_rsc_req_obj (
      .vd(din_0_rsc_req_obj_vd),
      .vz(din_0_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj_din_0_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj_din_0_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_0_rsc_req_obj_oswt(din_0_rsc_req_obj_oswt),
      .din_0_rsc_req_obj_vd(din_0_rsc_req_obj_vd),
      .din_0_rsc_req_obj_biwt(din_0_rsc_req_obj_biwt),
      .din_0_rsc_req_obj_bdwt(din_0_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj_din_0_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj_din_0_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_0_rsc_req_obj_oswt(din_0_rsc_req_obj_oswt),
      .din_0_rsc_req_obj_wen_comp(din_0_rsc_req_obj_wen_comp),
      .din_0_rsc_req_obj_biwt(din_0_rsc_req_obj_biwt),
      .din_0_rsc_req_obj_bdwt(din_0_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj (
  clk, rst, din_1_rsc_req_vz, core_wen, core_wten, din_1_rsc_req_obj_oswt, din_1_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_1_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_1_rsc_req_obj_oswt;
  output din_1_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_1_rsc_req_obj_vd;
  wire din_1_rsc_req_obj_biwt;
  wire din_1_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_1_rsc_req_obj (
      .vd(din_1_rsc_req_obj_vd),
      .vz(din_1_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj_din_1_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj_din_1_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_1_rsc_req_obj_oswt(din_1_rsc_req_obj_oswt),
      .din_1_rsc_req_obj_vd(din_1_rsc_req_obj_vd),
      .din_1_rsc_req_obj_biwt(din_1_rsc_req_obj_biwt),
      .din_1_rsc_req_obj_bdwt(din_1_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj_din_1_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj_din_1_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_1_rsc_req_obj_oswt(din_1_rsc_req_obj_oswt),
      .din_1_rsc_req_obj_wen_comp(din_1_rsc_req_obj_wen_comp),
      .din_1_rsc_req_obj_biwt(din_1_rsc_req_obj_biwt),
      .din_1_rsc_req_obj_bdwt(din_1_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj (
  clk, rst, din_2_rsc_req_vz, core_wen, core_wten, din_2_rsc_req_obj_oswt, din_2_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_2_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_2_rsc_req_obj_oswt;
  output din_2_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_2_rsc_req_obj_vd;
  wire din_2_rsc_req_obj_biwt;
  wire din_2_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_2_rsc_req_obj (
      .vd(din_2_rsc_req_obj_vd),
      .vz(din_2_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj_din_2_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj_din_2_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_2_rsc_req_obj_oswt(din_2_rsc_req_obj_oswt),
      .din_2_rsc_req_obj_vd(din_2_rsc_req_obj_vd),
      .din_2_rsc_req_obj_biwt(din_2_rsc_req_obj_biwt),
      .din_2_rsc_req_obj_bdwt(din_2_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj_din_2_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj_din_2_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_2_rsc_req_obj_oswt(din_2_rsc_req_obj_oswt),
      .din_2_rsc_req_obj_wen_comp(din_2_rsc_req_obj_wen_comp),
      .din_2_rsc_req_obj_biwt(din_2_rsc_req_obj_biwt),
      .din_2_rsc_req_obj_bdwt(din_2_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj (
  clk, rst, din_3_rsc_req_vz, core_wen, core_wten, din_3_rsc_req_obj_oswt, din_3_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_3_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_3_rsc_req_obj_oswt;
  output din_3_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_3_rsc_req_obj_vd;
  wire din_3_rsc_req_obj_biwt;
  wire din_3_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_3_rsc_req_obj (
      .vd(din_3_rsc_req_obj_vd),
      .vz(din_3_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj_din_3_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj_din_3_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_3_rsc_req_obj_oswt(din_3_rsc_req_obj_oswt),
      .din_3_rsc_req_obj_vd(din_3_rsc_req_obj_vd),
      .din_3_rsc_req_obj_biwt(din_3_rsc_req_obj_biwt),
      .din_3_rsc_req_obj_bdwt(din_3_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj_din_3_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj_din_3_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_3_rsc_req_obj_oswt(din_3_rsc_req_obj_oswt),
      .din_3_rsc_req_obj_wen_comp(din_3_rsc_req_obj_wen_comp),
      .din_3_rsc_req_obj_biwt(din_3_rsc_req_obj_biwt),
      .din_3_rsc_req_obj_bdwt(din_3_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj (
  clk, rst, din_4_rsc_req_vz, core_wen, core_wten, din_4_rsc_req_obj_oswt, din_4_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_4_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_4_rsc_req_obj_oswt;
  output din_4_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_4_rsc_req_obj_vd;
  wire din_4_rsc_req_obj_biwt;
  wire din_4_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_4_rsc_req_obj (
      .vd(din_4_rsc_req_obj_vd),
      .vz(din_4_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj_din_4_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj_din_4_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_4_rsc_req_obj_oswt(din_4_rsc_req_obj_oswt),
      .din_4_rsc_req_obj_vd(din_4_rsc_req_obj_vd),
      .din_4_rsc_req_obj_biwt(din_4_rsc_req_obj_biwt),
      .din_4_rsc_req_obj_bdwt(din_4_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj_din_4_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj_din_4_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_4_rsc_req_obj_oswt(din_4_rsc_req_obj_oswt),
      .din_4_rsc_req_obj_wen_comp(din_4_rsc_req_obj_wen_comp),
      .din_4_rsc_req_obj_biwt(din_4_rsc_req_obj_biwt),
      .din_4_rsc_req_obj_bdwt(din_4_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj (
  clk, rst, din_5_rsc_req_vz, core_wen, core_wten, din_5_rsc_req_obj_oswt, din_5_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_5_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_5_rsc_req_obj_oswt;
  output din_5_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_5_rsc_req_obj_vd;
  wire din_5_rsc_req_obj_biwt;
  wire din_5_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_5_rsc_req_obj (
      .vd(din_5_rsc_req_obj_vd),
      .vz(din_5_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj_din_5_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj_din_5_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_5_rsc_req_obj_oswt(din_5_rsc_req_obj_oswt),
      .din_5_rsc_req_obj_vd(din_5_rsc_req_obj_vd),
      .din_5_rsc_req_obj_biwt(din_5_rsc_req_obj_biwt),
      .din_5_rsc_req_obj_bdwt(din_5_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj_din_5_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj_din_5_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_5_rsc_req_obj_oswt(din_5_rsc_req_obj_oswt),
      .din_5_rsc_req_obj_wen_comp(din_5_rsc_req_obj_wen_comp),
      .din_5_rsc_req_obj_biwt(din_5_rsc_req_obj_biwt),
      .din_5_rsc_req_obj_bdwt(din_5_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj (
  clk, rst, din_6_rsc_req_vz, core_wen, core_wten, din_6_rsc_req_obj_oswt, din_6_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_6_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_6_rsc_req_obj_oswt;
  output din_6_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_6_rsc_req_obj_vd;
  wire din_6_rsc_req_obj_biwt;
  wire din_6_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_6_rsc_req_obj (
      .vd(din_6_rsc_req_obj_vd),
      .vz(din_6_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj_din_6_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj_din_6_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_6_rsc_req_obj_oswt(din_6_rsc_req_obj_oswt),
      .din_6_rsc_req_obj_vd(din_6_rsc_req_obj_vd),
      .din_6_rsc_req_obj_biwt(din_6_rsc_req_obj_biwt),
      .din_6_rsc_req_obj_bdwt(din_6_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj_din_6_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj_din_6_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_6_rsc_req_obj_oswt(din_6_rsc_req_obj_oswt),
      .din_6_rsc_req_obj_wen_comp(din_6_rsc_req_obj_wen_comp),
      .din_6_rsc_req_obj_biwt(din_6_rsc_req_obj_biwt),
      .din_6_rsc_req_obj_bdwt(din_6_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj (
  clk, rst, din_7_rsc_req_vz, core_wen, core_wten, din_7_rsc_req_obj_oswt, din_7_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_7_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_7_rsc_req_obj_oswt;
  output din_7_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_7_rsc_req_obj_vd;
  wire din_7_rsc_req_obj_biwt;
  wire din_7_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_7_rsc_req_obj (
      .vd(din_7_rsc_req_obj_vd),
      .vz(din_7_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj_din_7_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj_din_7_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_7_rsc_req_obj_oswt(din_7_rsc_req_obj_oswt),
      .din_7_rsc_req_obj_vd(din_7_rsc_req_obj_vd),
      .din_7_rsc_req_obj_biwt(din_7_rsc_req_obj_biwt),
      .din_7_rsc_req_obj_bdwt(din_7_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj_din_7_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj_din_7_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_7_rsc_req_obj_oswt(din_7_rsc_req_obj_oswt),
      .din_7_rsc_req_obj_wen_comp(din_7_rsc_req_obj_wen_comp),
      .din_7_rsc_req_obj_biwt(din_7_rsc_req_obj_biwt),
      .din_7_rsc_req_obj_bdwt(din_7_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj (
  clk, rst, din_8_rsc_req_vz, core_wen, core_wten, din_8_rsc_req_obj_oswt, din_8_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_8_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_8_rsc_req_obj_oswt;
  output din_8_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_8_rsc_req_obj_vd;
  wire din_8_rsc_req_obj_biwt;
  wire din_8_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_8_rsc_req_obj (
      .vd(din_8_rsc_req_obj_vd),
      .vz(din_8_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj_din_8_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj_din_8_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_8_rsc_req_obj_oswt(din_8_rsc_req_obj_oswt),
      .din_8_rsc_req_obj_vd(din_8_rsc_req_obj_vd),
      .din_8_rsc_req_obj_biwt(din_8_rsc_req_obj_biwt),
      .din_8_rsc_req_obj_bdwt(din_8_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj_din_8_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj_din_8_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_8_rsc_req_obj_oswt(din_8_rsc_req_obj_oswt),
      .din_8_rsc_req_obj_wen_comp(din_8_rsc_req_obj_wen_comp),
      .din_8_rsc_req_obj_biwt(din_8_rsc_req_obj_biwt),
      .din_8_rsc_req_obj_bdwt(din_8_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj (
  clk, rst, din_9_rsc_req_vz, core_wen, core_wten, din_9_rsc_req_obj_oswt, din_9_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_9_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_9_rsc_req_obj_oswt;
  output din_9_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_9_rsc_req_obj_vd;
  wire din_9_rsc_req_obj_biwt;
  wire din_9_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_9_rsc_req_obj (
      .vd(din_9_rsc_req_obj_vd),
      .vz(din_9_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj_din_9_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj_din_9_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_9_rsc_req_obj_oswt(din_9_rsc_req_obj_oswt),
      .din_9_rsc_req_obj_vd(din_9_rsc_req_obj_vd),
      .din_9_rsc_req_obj_biwt(din_9_rsc_req_obj_biwt),
      .din_9_rsc_req_obj_bdwt(din_9_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj_din_9_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj_din_9_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_9_rsc_req_obj_oswt(din_9_rsc_req_obj_oswt),
      .din_9_rsc_req_obj_wen_comp(din_9_rsc_req_obj_wen_comp),
      .din_9_rsc_req_obj_biwt(din_9_rsc_req_obj_biwt),
      .din_9_rsc_req_obj_bdwt(din_9_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj (
  clk, rst, din_10_rsc_req_vz, core_wen, core_wten, din_10_rsc_req_obj_oswt, din_10_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_10_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_10_rsc_req_obj_oswt;
  output din_10_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_10_rsc_req_obj_vd;
  wire din_10_rsc_req_obj_biwt;
  wire din_10_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_10_rsc_req_obj (
      .vd(din_10_rsc_req_obj_vd),
      .vz(din_10_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj_din_10_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj_din_10_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_10_rsc_req_obj_oswt(din_10_rsc_req_obj_oswt),
      .din_10_rsc_req_obj_vd(din_10_rsc_req_obj_vd),
      .din_10_rsc_req_obj_biwt(din_10_rsc_req_obj_biwt),
      .din_10_rsc_req_obj_bdwt(din_10_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj_din_10_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj_din_10_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_10_rsc_req_obj_oswt(din_10_rsc_req_obj_oswt),
      .din_10_rsc_req_obj_wen_comp(din_10_rsc_req_obj_wen_comp),
      .din_10_rsc_req_obj_biwt(din_10_rsc_req_obj_biwt),
      .din_10_rsc_req_obj_bdwt(din_10_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj (
  clk, rst, din_11_rsc_req_vz, core_wen, core_wten, din_11_rsc_req_obj_oswt, din_11_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_11_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_11_rsc_req_obj_oswt;
  output din_11_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_11_rsc_req_obj_vd;
  wire din_11_rsc_req_obj_biwt;
  wire din_11_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_11_rsc_req_obj (
      .vd(din_11_rsc_req_obj_vd),
      .vz(din_11_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj_din_11_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj_din_11_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_11_rsc_req_obj_oswt(din_11_rsc_req_obj_oswt),
      .din_11_rsc_req_obj_vd(din_11_rsc_req_obj_vd),
      .din_11_rsc_req_obj_biwt(din_11_rsc_req_obj_biwt),
      .din_11_rsc_req_obj_bdwt(din_11_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj_din_11_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj_din_11_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_11_rsc_req_obj_oswt(din_11_rsc_req_obj_oswt),
      .din_11_rsc_req_obj_wen_comp(din_11_rsc_req_obj_wen_comp),
      .din_11_rsc_req_obj_biwt(din_11_rsc_req_obj_biwt),
      .din_11_rsc_req_obj_bdwt(din_11_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj (
  clk, rst, din_12_rsc_req_vz, core_wen, core_wten, din_12_rsc_req_obj_oswt, din_12_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_12_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_12_rsc_req_obj_oswt;
  output din_12_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_12_rsc_req_obj_vd;
  wire din_12_rsc_req_obj_biwt;
  wire din_12_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_12_rsc_req_obj (
      .vd(din_12_rsc_req_obj_vd),
      .vz(din_12_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj_din_12_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj_din_12_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_12_rsc_req_obj_oswt(din_12_rsc_req_obj_oswt),
      .din_12_rsc_req_obj_vd(din_12_rsc_req_obj_vd),
      .din_12_rsc_req_obj_biwt(din_12_rsc_req_obj_biwt),
      .din_12_rsc_req_obj_bdwt(din_12_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj_din_12_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj_din_12_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_12_rsc_req_obj_oswt(din_12_rsc_req_obj_oswt),
      .din_12_rsc_req_obj_wen_comp(din_12_rsc_req_obj_wen_comp),
      .din_12_rsc_req_obj_biwt(din_12_rsc_req_obj_biwt),
      .din_12_rsc_req_obj_bdwt(din_12_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj (
  clk, rst, din_13_rsc_req_vz, core_wen, core_wten, din_13_rsc_req_obj_oswt, din_13_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_13_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_13_rsc_req_obj_oswt;
  output din_13_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_13_rsc_req_obj_vd;
  wire din_13_rsc_req_obj_biwt;
  wire din_13_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_13_rsc_req_obj (
      .vd(din_13_rsc_req_obj_vd),
      .vz(din_13_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj_din_13_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj_din_13_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_13_rsc_req_obj_oswt(din_13_rsc_req_obj_oswt),
      .din_13_rsc_req_obj_vd(din_13_rsc_req_obj_vd),
      .din_13_rsc_req_obj_biwt(din_13_rsc_req_obj_biwt),
      .din_13_rsc_req_obj_bdwt(din_13_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj_din_13_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj_din_13_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_13_rsc_req_obj_oswt(din_13_rsc_req_obj_oswt),
      .din_13_rsc_req_obj_wen_comp(din_13_rsc_req_obj_wen_comp),
      .din_13_rsc_req_obj_biwt(din_13_rsc_req_obj_biwt),
      .din_13_rsc_req_obj_bdwt(din_13_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj (
  clk, rst, din_14_rsc_req_vz, core_wen, core_wten, din_14_rsc_req_obj_oswt, din_14_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_14_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_14_rsc_req_obj_oswt;
  output din_14_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_14_rsc_req_obj_vd;
  wire din_14_rsc_req_obj_biwt;
  wire din_14_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_14_rsc_req_obj (
      .vd(din_14_rsc_req_obj_vd),
      .vz(din_14_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj_din_14_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj_din_14_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_14_rsc_req_obj_oswt(din_14_rsc_req_obj_oswt),
      .din_14_rsc_req_obj_vd(din_14_rsc_req_obj_vd),
      .din_14_rsc_req_obj_biwt(din_14_rsc_req_obj_biwt),
      .din_14_rsc_req_obj_bdwt(din_14_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj_din_14_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj_din_14_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_14_rsc_req_obj_oswt(din_14_rsc_req_obj_oswt),
      .din_14_rsc_req_obj_wen_comp(din_14_rsc_req_obj_wen_comp),
      .din_14_rsc_req_obj_biwt(din_14_rsc_req_obj_biwt),
      .din_14_rsc_req_obj_bdwt(din_14_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj (
  clk, rst, din_15_rsc_req_vz, core_wen, core_wten, din_15_rsc_req_obj_oswt, din_15_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_15_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_15_rsc_req_obj_oswt;
  output din_15_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_15_rsc_req_obj_vd;
  wire din_15_rsc_req_obj_biwt;
  wire din_15_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_15_rsc_req_obj (
      .vd(din_15_rsc_req_obj_vd),
      .vz(din_15_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj_din_15_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj_din_15_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_15_rsc_req_obj_oswt(din_15_rsc_req_obj_oswt),
      .din_15_rsc_req_obj_vd(din_15_rsc_req_obj_vd),
      .din_15_rsc_req_obj_biwt(din_15_rsc_req_obj_biwt),
      .din_15_rsc_req_obj_bdwt(din_15_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj_din_15_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj_din_15_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_15_rsc_req_obj_oswt(din_15_rsc_req_obj_oswt),
      .din_15_rsc_req_obj_wen_comp(din_15_rsc_req_obj_wen_comp),
      .din_15_rsc_req_obj_biwt(din_15_rsc_req_obj_biwt),
      .din_15_rsc_req_obj_bdwt(din_15_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj (
  clk, rst, din_16_rsc_req_vz, core_wen, core_wten, din_16_rsc_req_obj_oswt, din_16_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_16_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_16_rsc_req_obj_oswt;
  output din_16_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_16_rsc_req_obj_vd;
  wire din_16_rsc_req_obj_biwt;
  wire din_16_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_16_rsc_req_obj (
      .vd(din_16_rsc_req_obj_vd),
      .vz(din_16_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj_din_16_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj_din_16_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_16_rsc_req_obj_oswt(din_16_rsc_req_obj_oswt),
      .din_16_rsc_req_obj_vd(din_16_rsc_req_obj_vd),
      .din_16_rsc_req_obj_biwt(din_16_rsc_req_obj_biwt),
      .din_16_rsc_req_obj_bdwt(din_16_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj_din_16_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj_din_16_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_16_rsc_req_obj_oswt(din_16_rsc_req_obj_oswt),
      .din_16_rsc_req_obj_wen_comp(din_16_rsc_req_obj_wen_comp),
      .din_16_rsc_req_obj_biwt(din_16_rsc_req_obj_biwt),
      .din_16_rsc_req_obj_bdwt(din_16_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj (
  clk, rst, din_17_rsc_req_vz, core_wen, core_wten, din_17_rsc_req_obj_oswt, din_17_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_17_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_17_rsc_req_obj_oswt;
  output din_17_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_17_rsc_req_obj_vd;
  wire din_17_rsc_req_obj_biwt;
  wire din_17_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_17_rsc_req_obj (
      .vd(din_17_rsc_req_obj_vd),
      .vz(din_17_rsc_req_vz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj_din_17_rsc_req_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj_din_17_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_17_rsc_req_obj_oswt(din_17_rsc_req_obj_oswt),
      .din_17_rsc_req_obj_vd(din_17_rsc_req_obj_vd),
      .din_17_rsc_req_obj_biwt(din_17_rsc_req_obj_biwt),
      .din_17_rsc_req_obj_bdwt(din_17_rsc_req_obj_bdwt)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj_din_17_rsc_req_wait_dp
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj_din_17_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_17_rsc_req_obj_oswt(din_17_rsc_req_obj_oswt),
      .din_17_rsc_req_obj_wen_comp(din_17_rsc_req_obj_wen_comp),
      .din_17_rsc_req_obj_biwt(din_17_rsc_req_obj_biwt),
      .din_17_rsc_req_obj_bdwt(din_17_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_rls_obj (
  din_17_rsc_rls_lz, core_wten, din_17_rsc_rls_obj_iswt0
);
  output din_17_rsc_rls_lz;
  input core_wten;
  input din_17_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_17_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_17_rsc_rls_obj (
      .ld(din_17_rsc_rls_obj_ld_core_sct),
      .lz(din_17_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_rls_obj_din_17_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_rls_obj_din_17_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_17_rsc_rls_obj_iswt0(din_17_rsc_rls_obj_iswt0),
      .din_17_rsc_rls_obj_ld_core_sct(din_17_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_rls_obj (
  din_16_rsc_rls_lz, core_wten, din_16_rsc_rls_obj_iswt0
);
  output din_16_rsc_rls_lz;
  input core_wten;
  input din_16_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_16_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_16_rsc_rls_obj (
      .ld(din_16_rsc_rls_obj_ld_core_sct),
      .lz(din_16_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_rls_obj_din_16_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_rls_obj_din_16_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_16_rsc_rls_obj_iswt0(din_16_rsc_rls_obj_iswt0),
      .din_16_rsc_rls_obj_ld_core_sct(din_16_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_rls_obj (
  din_15_rsc_rls_lz, core_wten, din_15_rsc_rls_obj_iswt0
);
  output din_15_rsc_rls_lz;
  input core_wten;
  input din_15_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_15_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_15_rsc_rls_obj (
      .ld(din_15_rsc_rls_obj_ld_core_sct),
      .lz(din_15_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_rls_obj_din_15_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_rls_obj_din_15_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_15_rsc_rls_obj_iswt0(din_15_rsc_rls_obj_iswt0),
      .din_15_rsc_rls_obj_ld_core_sct(din_15_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_rls_obj (
  din_14_rsc_rls_lz, core_wten, din_14_rsc_rls_obj_iswt0
);
  output din_14_rsc_rls_lz;
  input core_wten;
  input din_14_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_14_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_14_rsc_rls_obj (
      .ld(din_14_rsc_rls_obj_ld_core_sct),
      .lz(din_14_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_rls_obj_din_14_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_rls_obj_din_14_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_14_rsc_rls_obj_iswt0(din_14_rsc_rls_obj_iswt0),
      .din_14_rsc_rls_obj_ld_core_sct(din_14_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_rls_obj (
  din_13_rsc_rls_lz, core_wten, din_13_rsc_rls_obj_iswt0
);
  output din_13_rsc_rls_lz;
  input core_wten;
  input din_13_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_13_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_13_rsc_rls_obj (
      .ld(din_13_rsc_rls_obj_ld_core_sct),
      .lz(din_13_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_rls_obj_din_13_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_rls_obj_din_13_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_13_rsc_rls_obj_iswt0(din_13_rsc_rls_obj_iswt0),
      .din_13_rsc_rls_obj_ld_core_sct(din_13_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_rls_obj (
  din_12_rsc_rls_lz, core_wten, din_12_rsc_rls_obj_iswt0
);
  output din_12_rsc_rls_lz;
  input core_wten;
  input din_12_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_12_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_12_rsc_rls_obj (
      .ld(din_12_rsc_rls_obj_ld_core_sct),
      .lz(din_12_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_rls_obj_din_12_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_rls_obj_din_12_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_12_rsc_rls_obj_iswt0(din_12_rsc_rls_obj_iswt0),
      .din_12_rsc_rls_obj_ld_core_sct(din_12_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_rls_obj (
  din_11_rsc_rls_lz, core_wten, din_11_rsc_rls_obj_iswt0
);
  output din_11_rsc_rls_lz;
  input core_wten;
  input din_11_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_11_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_11_rsc_rls_obj (
      .ld(din_11_rsc_rls_obj_ld_core_sct),
      .lz(din_11_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_rls_obj_din_11_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_rls_obj_din_11_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_11_rsc_rls_obj_iswt0(din_11_rsc_rls_obj_iswt0),
      .din_11_rsc_rls_obj_ld_core_sct(din_11_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_rls_obj (
  din_10_rsc_rls_lz, core_wten, din_10_rsc_rls_obj_iswt0
);
  output din_10_rsc_rls_lz;
  input core_wten;
  input din_10_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_10_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_10_rsc_rls_obj (
      .ld(din_10_rsc_rls_obj_ld_core_sct),
      .lz(din_10_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_rls_obj_din_10_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_rls_obj_din_10_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_10_rsc_rls_obj_iswt0(din_10_rsc_rls_obj_iswt0),
      .din_10_rsc_rls_obj_ld_core_sct(din_10_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_rls_obj (
  din_9_rsc_rls_lz, core_wten, din_9_rsc_rls_obj_iswt0
);
  output din_9_rsc_rls_lz;
  input core_wten;
  input din_9_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_9_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_9_rsc_rls_obj (
      .ld(din_9_rsc_rls_obj_ld_core_sct),
      .lz(din_9_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_rls_obj_din_9_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_rls_obj_din_9_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_9_rsc_rls_obj_iswt0(din_9_rsc_rls_obj_iswt0),
      .din_9_rsc_rls_obj_ld_core_sct(din_9_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_rls_obj (
  din_8_rsc_rls_lz, core_wten, din_8_rsc_rls_obj_iswt0
);
  output din_8_rsc_rls_lz;
  input core_wten;
  input din_8_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_8_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_8_rsc_rls_obj (
      .ld(din_8_rsc_rls_obj_ld_core_sct),
      .lz(din_8_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_rls_obj_din_8_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_rls_obj_din_8_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_8_rsc_rls_obj_iswt0(din_8_rsc_rls_obj_iswt0),
      .din_8_rsc_rls_obj_ld_core_sct(din_8_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_rls_obj (
  din_7_rsc_rls_lz, core_wten, din_7_rsc_rls_obj_iswt0
);
  output din_7_rsc_rls_lz;
  input core_wten;
  input din_7_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_7_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_7_rsc_rls_obj (
      .ld(din_7_rsc_rls_obj_ld_core_sct),
      .lz(din_7_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_rls_obj_din_7_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_rls_obj_din_7_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_7_rsc_rls_obj_iswt0(din_7_rsc_rls_obj_iswt0),
      .din_7_rsc_rls_obj_ld_core_sct(din_7_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_rls_obj (
  din_6_rsc_rls_lz, core_wten, din_6_rsc_rls_obj_iswt0
);
  output din_6_rsc_rls_lz;
  input core_wten;
  input din_6_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_6_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_6_rsc_rls_obj (
      .ld(din_6_rsc_rls_obj_ld_core_sct),
      .lz(din_6_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_rls_obj_din_6_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_rls_obj_din_6_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_6_rsc_rls_obj_iswt0(din_6_rsc_rls_obj_iswt0),
      .din_6_rsc_rls_obj_ld_core_sct(din_6_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_rls_obj (
  din_5_rsc_rls_lz, core_wten, din_5_rsc_rls_obj_iswt0
);
  output din_5_rsc_rls_lz;
  input core_wten;
  input din_5_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_5_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_5_rsc_rls_obj (
      .ld(din_5_rsc_rls_obj_ld_core_sct),
      .lz(din_5_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_rls_obj_din_5_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_rls_obj_din_5_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_5_rsc_rls_obj_iswt0(din_5_rsc_rls_obj_iswt0),
      .din_5_rsc_rls_obj_ld_core_sct(din_5_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_rls_obj (
  din_4_rsc_rls_lz, core_wten, din_4_rsc_rls_obj_iswt0
);
  output din_4_rsc_rls_lz;
  input core_wten;
  input din_4_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_4_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_4_rsc_rls_obj (
      .ld(din_4_rsc_rls_obj_ld_core_sct),
      .lz(din_4_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_rls_obj_din_4_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_rls_obj_din_4_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_4_rsc_rls_obj_iswt0(din_4_rsc_rls_obj_iswt0),
      .din_4_rsc_rls_obj_ld_core_sct(din_4_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_rls_obj (
  din_3_rsc_rls_lz, core_wten, din_3_rsc_rls_obj_iswt0
);
  output din_3_rsc_rls_lz;
  input core_wten;
  input din_3_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_3_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_3_rsc_rls_obj (
      .ld(din_3_rsc_rls_obj_ld_core_sct),
      .lz(din_3_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_rls_obj_din_3_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_rls_obj_din_3_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_3_rsc_rls_obj_iswt0(din_3_rsc_rls_obj_iswt0),
      .din_3_rsc_rls_obj_ld_core_sct(din_3_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_rls_obj (
  din_2_rsc_rls_lz, core_wten, din_2_rsc_rls_obj_iswt0
);
  output din_2_rsc_rls_lz;
  input core_wten;
  input din_2_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_2_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_2_rsc_rls_obj (
      .ld(din_2_rsc_rls_obj_ld_core_sct),
      .lz(din_2_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_rls_obj_din_2_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_rls_obj_din_2_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_2_rsc_rls_obj_iswt0(din_2_rsc_rls_obj_iswt0),
      .din_2_rsc_rls_obj_ld_core_sct(din_2_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_rls_obj (
  din_1_rsc_rls_lz, core_wten, din_1_rsc_rls_obj_iswt0
);
  output din_1_rsc_rls_lz;
  input core_wten;
  input din_1_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_1_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_1_rsc_rls_obj (
      .ld(din_1_rsc_rls_obj_ld_core_sct),
      .lz(din_1_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_rls_obj_din_1_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_rls_obj_din_1_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_1_rsc_rls_obj_iswt0(din_1_rsc_rls_obj_iswt0),
      .din_1_rsc_rls_obj_ld_core_sct(din_1_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_rls_obj (
  din_0_rsc_rls_lz, core_wten, din_0_rsc_rls_obj_iswt0
);
  output din_0_rsc_rls_lz;
  input core_wten;
  input din_0_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_0_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_0_rsc_rls_obj (
      .ld(din_0_rsc_rls_obj_ld_core_sct),
      .lz(din_0_rsc_rls_lz)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_rls_obj_din_0_rsc_rls_wait_ctrl
      READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_rls_obj_din_0_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_0_rsc_rls_obj_iswt0(din_0_rsc_rls_obj_iswt0),
      .din_0_rsc_rls_obj_ld_core_sct(din_0_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci (
  clk, rst, dout_rsc_z, dout_rsc_vz, dout_rsc_lz, core_wen, core_wten, dout_rsci_oswt,
      dout_rsci_wen_comp, dout_rsci_d
);
  input clk;
  input rst;
  output [511:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;
  input core_wen;
  input core_wten;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input [511:0] dout_rsci_d;


  // Interconnect Declarations
  wire dout_rsci_biwt;
  wire dout_rsci_bdwt;
  wire dout_rsci_ld_core_sct;
  wire dout_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  mgc_out_stdreg_wait_v1 #(.rscid(32'sd56),
  .width(32'sd512)) dout_rsci (
      .ld(dout_rsci_ld_core_sct),
      .vd(dout_rsci_vd),
      .d(dout_rsci_d),
      .lz(dout_rsc_lz),
      .vz(dout_rsc_vz),
      .z(dout_rsc_z)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_dout_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_dout_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_ld_core_sct(dout_rsci_ld_core_sct),
      .dout_rsci_vd(dout_rsci_vd)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_dout_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_dout_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1 (
  clk, rst, din_17_rsci_douta_d, din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_17_rsci_oswt, din_17_rsci_douta_d_mxwt, din_17_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_17_rsci_douta_d;
  output din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_17_rsci_oswt;
  output [15:0] din_17_rsci_douta_d_mxwt;
  input din_17_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_17_rsci_biwt;
  wire din_17_rsci_bdwt;
  wire [15:0] din_17_rsci_douta_d_mxwt_pconst;
  wire din_17_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1_din_17_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1_din_17_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_17_rsci_oswt(din_17_rsci_oswt),
      .din_17_rsci_biwt(din_17_rsci_biwt),
      .din_17_rsci_bdwt(din_17_rsci_bdwt),
      .din_17_rsci_biwt_pff(din_17_rsci_biwt_iff),
      .din_17_rsci_oswt_pff(din_17_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1_din_17_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1_din_17_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_17_rsci_douta_d(din_17_rsci_douta_d),
      .din_17_rsci_douta_d_mxwt(din_17_rsci_douta_d_mxwt_pconst),
      .din_17_rsci_biwt(din_17_rsci_biwt),
      .din_17_rsci_bdwt(din_17_rsci_bdwt)
    );
  assign din_17_rsci_douta_d_mxwt = din_17_rsci_douta_d_mxwt_pconst;
  assign din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_17_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1 (
  clk, rst, din_16_rsci_douta_d, din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_16_rsci_oswt, din_16_rsci_douta_d_mxwt, din_16_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_16_rsci_douta_d;
  output din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_16_rsci_oswt;
  output [15:0] din_16_rsci_douta_d_mxwt;
  input din_16_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_16_rsci_biwt;
  wire din_16_rsci_bdwt;
  wire [15:0] din_16_rsci_douta_d_mxwt_pconst;
  wire din_16_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1_din_16_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1_din_16_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_16_rsci_oswt(din_16_rsci_oswt),
      .din_16_rsci_biwt(din_16_rsci_biwt),
      .din_16_rsci_bdwt(din_16_rsci_bdwt),
      .din_16_rsci_biwt_pff(din_16_rsci_biwt_iff),
      .din_16_rsci_oswt_pff(din_16_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1_din_16_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1_din_16_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_16_rsci_douta_d(din_16_rsci_douta_d),
      .din_16_rsci_douta_d_mxwt(din_16_rsci_douta_d_mxwt_pconst),
      .din_16_rsci_biwt(din_16_rsci_biwt),
      .din_16_rsci_bdwt(din_16_rsci_bdwt)
    );
  assign din_16_rsci_douta_d_mxwt = din_16_rsci_douta_d_mxwt_pconst;
  assign din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_16_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1 (
  clk, rst, din_15_rsci_douta_d, din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_15_rsci_oswt, din_15_rsci_douta_d_mxwt, din_15_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_15_rsci_douta_d;
  output din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_15_rsci_oswt;
  output [15:0] din_15_rsci_douta_d_mxwt;
  input din_15_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_15_rsci_biwt;
  wire din_15_rsci_bdwt;
  wire [15:0] din_15_rsci_douta_d_mxwt_pconst;
  wire din_15_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1_din_15_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1_din_15_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_15_rsci_oswt(din_15_rsci_oswt),
      .din_15_rsci_biwt(din_15_rsci_biwt),
      .din_15_rsci_bdwt(din_15_rsci_bdwt),
      .din_15_rsci_biwt_pff(din_15_rsci_biwt_iff),
      .din_15_rsci_oswt_pff(din_15_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1_din_15_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1_din_15_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_15_rsci_douta_d(din_15_rsci_douta_d),
      .din_15_rsci_douta_d_mxwt(din_15_rsci_douta_d_mxwt_pconst),
      .din_15_rsci_biwt(din_15_rsci_biwt),
      .din_15_rsci_bdwt(din_15_rsci_bdwt)
    );
  assign din_15_rsci_douta_d_mxwt = din_15_rsci_douta_d_mxwt_pconst;
  assign din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_15_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1 (
  clk, rst, din_14_rsci_douta_d, din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_14_rsci_oswt, din_14_rsci_douta_d_mxwt, din_14_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_14_rsci_douta_d;
  output din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_14_rsci_oswt;
  output [15:0] din_14_rsci_douta_d_mxwt;
  input din_14_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_14_rsci_biwt;
  wire din_14_rsci_bdwt;
  wire [15:0] din_14_rsci_douta_d_mxwt_pconst;
  wire din_14_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1_din_14_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1_din_14_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_14_rsci_oswt(din_14_rsci_oswt),
      .din_14_rsci_biwt(din_14_rsci_biwt),
      .din_14_rsci_bdwt(din_14_rsci_bdwt),
      .din_14_rsci_biwt_pff(din_14_rsci_biwt_iff),
      .din_14_rsci_oswt_pff(din_14_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1_din_14_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1_din_14_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_14_rsci_douta_d(din_14_rsci_douta_d),
      .din_14_rsci_douta_d_mxwt(din_14_rsci_douta_d_mxwt_pconst),
      .din_14_rsci_biwt(din_14_rsci_biwt),
      .din_14_rsci_bdwt(din_14_rsci_bdwt)
    );
  assign din_14_rsci_douta_d_mxwt = din_14_rsci_douta_d_mxwt_pconst;
  assign din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_14_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1 (
  clk, rst, din_13_rsci_douta_d, din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_13_rsci_oswt, din_13_rsci_douta_d_mxwt, din_13_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_13_rsci_douta_d;
  output din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_13_rsci_oswt;
  output [15:0] din_13_rsci_douta_d_mxwt;
  input din_13_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_13_rsci_biwt;
  wire din_13_rsci_bdwt;
  wire [15:0] din_13_rsci_douta_d_mxwt_pconst;
  wire din_13_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1_din_13_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1_din_13_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_13_rsci_oswt(din_13_rsci_oswt),
      .din_13_rsci_biwt(din_13_rsci_biwt),
      .din_13_rsci_bdwt(din_13_rsci_bdwt),
      .din_13_rsci_biwt_pff(din_13_rsci_biwt_iff),
      .din_13_rsci_oswt_pff(din_13_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1_din_13_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1_din_13_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_13_rsci_douta_d(din_13_rsci_douta_d),
      .din_13_rsci_douta_d_mxwt(din_13_rsci_douta_d_mxwt_pconst),
      .din_13_rsci_biwt(din_13_rsci_biwt),
      .din_13_rsci_bdwt(din_13_rsci_bdwt)
    );
  assign din_13_rsci_douta_d_mxwt = din_13_rsci_douta_d_mxwt_pconst;
  assign din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_13_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1 (
  clk, rst, din_12_rsci_douta_d, din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_12_rsci_oswt, din_12_rsci_douta_d_mxwt, din_12_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_12_rsci_douta_d;
  output din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_12_rsci_oswt;
  output [15:0] din_12_rsci_douta_d_mxwt;
  input din_12_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_12_rsci_biwt;
  wire din_12_rsci_bdwt;
  wire [15:0] din_12_rsci_douta_d_mxwt_pconst;
  wire din_12_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1_din_12_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1_din_12_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_12_rsci_oswt(din_12_rsci_oswt),
      .din_12_rsci_biwt(din_12_rsci_biwt),
      .din_12_rsci_bdwt(din_12_rsci_bdwt),
      .din_12_rsci_biwt_pff(din_12_rsci_biwt_iff),
      .din_12_rsci_oswt_pff(din_12_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1_din_12_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1_din_12_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_12_rsci_douta_d(din_12_rsci_douta_d),
      .din_12_rsci_douta_d_mxwt(din_12_rsci_douta_d_mxwt_pconst),
      .din_12_rsci_biwt(din_12_rsci_biwt),
      .din_12_rsci_bdwt(din_12_rsci_bdwt)
    );
  assign din_12_rsci_douta_d_mxwt = din_12_rsci_douta_d_mxwt_pconst;
  assign din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_12_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1 (
  clk, rst, din_11_rsci_douta_d, din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_11_rsci_oswt, din_11_rsci_douta_d_mxwt, din_11_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_11_rsci_douta_d;
  output din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_11_rsci_oswt;
  output [15:0] din_11_rsci_douta_d_mxwt;
  input din_11_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_11_rsci_biwt;
  wire din_11_rsci_bdwt;
  wire [15:0] din_11_rsci_douta_d_mxwt_pconst;
  wire din_11_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1_din_11_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1_din_11_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_11_rsci_oswt(din_11_rsci_oswt),
      .din_11_rsci_biwt(din_11_rsci_biwt),
      .din_11_rsci_bdwt(din_11_rsci_bdwt),
      .din_11_rsci_biwt_pff(din_11_rsci_biwt_iff),
      .din_11_rsci_oswt_pff(din_11_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1_din_11_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1_din_11_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_11_rsci_douta_d(din_11_rsci_douta_d),
      .din_11_rsci_douta_d_mxwt(din_11_rsci_douta_d_mxwt_pconst),
      .din_11_rsci_biwt(din_11_rsci_biwt),
      .din_11_rsci_bdwt(din_11_rsci_bdwt)
    );
  assign din_11_rsci_douta_d_mxwt = din_11_rsci_douta_d_mxwt_pconst;
  assign din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_11_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1 (
  clk, rst, din_10_rsci_douta_d, din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_10_rsci_oswt, din_10_rsci_douta_d_mxwt, din_10_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_10_rsci_douta_d;
  output din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_10_rsci_oswt;
  output [15:0] din_10_rsci_douta_d_mxwt;
  input din_10_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_10_rsci_biwt;
  wire din_10_rsci_bdwt;
  wire [15:0] din_10_rsci_douta_d_mxwt_pconst;
  wire din_10_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1_din_10_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1_din_10_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_10_rsci_oswt(din_10_rsci_oswt),
      .din_10_rsci_biwt(din_10_rsci_biwt),
      .din_10_rsci_bdwt(din_10_rsci_bdwt),
      .din_10_rsci_biwt_pff(din_10_rsci_biwt_iff),
      .din_10_rsci_oswt_pff(din_10_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1_din_10_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1_din_10_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_10_rsci_douta_d(din_10_rsci_douta_d),
      .din_10_rsci_douta_d_mxwt(din_10_rsci_douta_d_mxwt_pconst),
      .din_10_rsci_biwt(din_10_rsci_biwt),
      .din_10_rsci_bdwt(din_10_rsci_bdwt)
    );
  assign din_10_rsci_douta_d_mxwt = din_10_rsci_douta_d_mxwt_pconst;
  assign din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_10_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1 (
  clk, rst, din_9_rsci_douta_d, din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_9_rsci_oswt, din_9_rsci_douta_d_mxwt, din_9_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_9_rsci_douta_d;
  output din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_9_rsci_oswt;
  output [15:0] din_9_rsci_douta_d_mxwt;
  input din_9_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_9_rsci_biwt;
  wire din_9_rsci_bdwt;
  wire [15:0] din_9_rsci_douta_d_mxwt_pconst;
  wire din_9_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1_din_9_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1_din_9_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_9_rsci_oswt(din_9_rsci_oswt),
      .din_9_rsci_biwt(din_9_rsci_biwt),
      .din_9_rsci_bdwt(din_9_rsci_bdwt),
      .din_9_rsci_biwt_pff(din_9_rsci_biwt_iff),
      .din_9_rsci_oswt_pff(din_9_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1_din_9_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1_din_9_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_9_rsci_douta_d(din_9_rsci_douta_d),
      .din_9_rsci_douta_d_mxwt(din_9_rsci_douta_d_mxwt_pconst),
      .din_9_rsci_biwt(din_9_rsci_biwt),
      .din_9_rsci_bdwt(din_9_rsci_bdwt)
    );
  assign din_9_rsci_douta_d_mxwt = din_9_rsci_douta_d_mxwt_pconst;
  assign din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_9_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1 (
  clk, rst, din_8_rsci_douta_d, din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_8_rsci_oswt, din_8_rsci_douta_d_mxwt, din_8_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_8_rsci_douta_d;
  output din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_8_rsci_oswt;
  output [15:0] din_8_rsci_douta_d_mxwt;
  input din_8_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_8_rsci_biwt;
  wire din_8_rsci_bdwt;
  wire [15:0] din_8_rsci_douta_d_mxwt_pconst;
  wire din_8_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1_din_8_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1_din_8_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_8_rsci_oswt(din_8_rsci_oswt),
      .din_8_rsci_biwt(din_8_rsci_biwt),
      .din_8_rsci_bdwt(din_8_rsci_bdwt),
      .din_8_rsci_biwt_pff(din_8_rsci_biwt_iff),
      .din_8_rsci_oswt_pff(din_8_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1_din_8_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1_din_8_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_8_rsci_douta_d(din_8_rsci_douta_d),
      .din_8_rsci_douta_d_mxwt(din_8_rsci_douta_d_mxwt_pconst),
      .din_8_rsci_biwt(din_8_rsci_biwt),
      .din_8_rsci_bdwt(din_8_rsci_bdwt)
    );
  assign din_8_rsci_douta_d_mxwt = din_8_rsci_douta_d_mxwt_pconst;
  assign din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_8_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1 (
  clk, rst, din_7_rsci_douta_d, din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_7_rsci_oswt, din_7_rsci_douta_d_mxwt, din_7_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_7_rsci_douta_d;
  output din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_7_rsci_oswt;
  output [15:0] din_7_rsci_douta_d_mxwt;
  input din_7_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_7_rsci_biwt;
  wire din_7_rsci_bdwt;
  wire [15:0] din_7_rsci_douta_d_mxwt_pconst;
  wire din_7_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1_din_7_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1_din_7_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_7_rsci_oswt(din_7_rsci_oswt),
      .din_7_rsci_biwt(din_7_rsci_biwt),
      .din_7_rsci_bdwt(din_7_rsci_bdwt),
      .din_7_rsci_biwt_pff(din_7_rsci_biwt_iff),
      .din_7_rsci_oswt_pff(din_7_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1_din_7_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1_din_7_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_7_rsci_douta_d(din_7_rsci_douta_d),
      .din_7_rsci_douta_d_mxwt(din_7_rsci_douta_d_mxwt_pconst),
      .din_7_rsci_biwt(din_7_rsci_biwt),
      .din_7_rsci_bdwt(din_7_rsci_bdwt)
    );
  assign din_7_rsci_douta_d_mxwt = din_7_rsci_douta_d_mxwt_pconst;
  assign din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_7_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1 (
  clk, rst, din_6_rsci_douta_d, din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_6_rsci_oswt, din_6_rsci_douta_d_mxwt, din_6_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_6_rsci_douta_d;
  output din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_6_rsci_oswt;
  output [15:0] din_6_rsci_douta_d_mxwt;
  input din_6_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_6_rsci_biwt;
  wire din_6_rsci_bdwt;
  wire [15:0] din_6_rsci_douta_d_mxwt_pconst;
  wire din_6_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1_din_6_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1_din_6_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_6_rsci_oswt(din_6_rsci_oswt),
      .din_6_rsci_biwt(din_6_rsci_biwt),
      .din_6_rsci_bdwt(din_6_rsci_bdwt),
      .din_6_rsci_biwt_pff(din_6_rsci_biwt_iff),
      .din_6_rsci_oswt_pff(din_6_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1_din_6_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1_din_6_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_6_rsci_douta_d(din_6_rsci_douta_d),
      .din_6_rsci_douta_d_mxwt(din_6_rsci_douta_d_mxwt_pconst),
      .din_6_rsci_biwt(din_6_rsci_biwt),
      .din_6_rsci_bdwt(din_6_rsci_bdwt)
    );
  assign din_6_rsci_douta_d_mxwt = din_6_rsci_douta_d_mxwt_pconst;
  assign din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_6_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1 (
  clk, rst, din_5_rsci_douta_d, din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_5_rsci_oswt, din_5_rsci_douta_d_mxwt, din_5_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_5_rsci_douta_d;
  output din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_5_rsci_oswt;
  output [15:0] din_5_rsci_douta_d_mxwt;
  input din_5_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_5_rsci_biwt;
  wire din_5_rsci_bdwt;
  wire [15:0] din_5_rsci_douta_d_mxwt_pconst;
  wire din_5_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1_din_5_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1_din_5_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_5_rsci_oswt(din_5_rsci_oswt),
      .din_5_rsci_biwt(din_5_rsci_biwt),
      .din_5_rsci_bdwt(din_5_rsci_bdwt),
      .din_5_rsci_biwt_pff(din_5_rsci_biwt_iff),
      .din_5_rsci_oswt_pff(din_5_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1_din_5_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1_din_5_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_5_rsci_douta_d(din_5_rsci_douta_d),
      .din_5_rsci_douta_d_mxwt(din_5_rsci_douta_d_mxwt_pconst),
      .din_5_rsci_biwt(din_5_rsci_biwt),
      .din_5_rsci_bdwt(din_5_rsci_bdwt)
    );
  assign din_5_rsci_douta_d_mxwt = din_5_rsci_douta_d_mxwt_pconst;
  assign din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_5_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1 (
  clk, rst, din_4_rsci_douta_d, din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_4_rsci_oswt, din_4_rsci_douta_d_mxwt, din_4_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_4_rsci_douta_d;
  output din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_4_rsci_oswt;
  output [15:0] din_4_rsci_douta_d_mxwt;
  input din_4_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_4_rsci_biwt;
  wire din_4_rsci_bdwt;
  wire [15:0] din_4_rsci_douta_d_mxwt_pconst;
  wire din_4_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1_din_4_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1_din_4_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_4_rsci_oswt(din_4_rsci_oswt),
      .din_4_rsci_biwt(din_4_rsci_biwt),
      .din_4_rsci_bdwt(din_4_rsci_bdwt),
      .din_4_rsci_biwt_pff(din_4_rsci_biwt_iff),
      .din_4_rsci_oswt_pff(din_4_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1_din_4_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1_din_4_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_4_rsci_douta_d(din_4_rsci_douta_d),
      .din_4_rsci_douta_d_mxwt(din_4_rsci_douta_d_mxwt_pconst),
      .din_4_rsci_biwt(din_4_rsci_biwt),
      .din_4_rsci_bdwt(din_4_rsci_bdwt)
    );
  assign din_4_rsci_douta_d_mxwt = din_4_rsci_douta_d_mxwt_pconst;
  assign din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_4_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1 (
  clk, rst, din_3_rsci_douta_d, din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_3_rsci_oswt, din_3_rsci_douta_d_mxwt, din_3_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_3_rsci_douta_d;
  output din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_3_rsci_oswt;
  output [15:0] din_3_rsci_douta_d_mxwt;
  input din_3_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_3_rsci_biwt;
  wire din_3_rsci_bdwt;
  wire [15:0] din_3_rsci_douta_d_mxwt_pconst;
  wire din_3_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1_din_3_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1_din_3_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_3_rsci_oswt(din_3_rsci_oswt),
      .din_3_rsci_biwt(din_3_rsci_biwt),
      .din_3_rsci_bdwt(din_3_rsci_bdwt),
      .din_3_rsci_biwt_pff(din_3_rsci_biwt_iff),
      .din_3_rsci_oswt_pff(din_3_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1_din_3_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1_din_3_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_3_rsci_douta_d(din_3_rsci_douta_d),
      .din_3_rsci_douta_d_mxwt(din_3_rsci_douta_d_mxwt_pconst),
      .din_3_rsci_biwt(din_3_rsci_biwt),
      .din_3_rsci_bdwt(din_3_rsci_bdwt)
    );
  assign din_3_rsci_douta_d_mxwt = din_3_rsci_douta_d_mxwt_pconst;
  assign din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_3_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1 (
  clk, rst, din_2_rsci_douta_d, din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_2_rsci_oswt, din_2_rsci_douta_d_mxwt, din_2_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_2_rsci_douta_d;
  output din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_2_rsci_oswt;
  output [15:0] din_2_rsci_douta_d_mxwt;
  input din_2_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_2_rsci_biwt;
  wire din_2_rsci_bdwt;
  wire [15:0] din_2_rsci_douta_d_mxwt_pconst;
  wire din_2_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1_din_2_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1_din_2_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_2_rsci_oswt(din_2_rsci_oswt),
      .din_2_rsci_biwt(din_2_rsci_biwt),
      .din_2_rsci_bdwt(din_2_rsci_bdwt),
      .din_2_rsci_biwt_pff(din_2_rsci_biwt_iff),
      .din_2_rsci_oswt_pff(din_2_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1_din_2_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1_din_2_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_2_rsci_douta_d(din_2_rsci_douta_d),
      .din_2_rsci_douta_d_mxwt(din_2_rsci_douta_d_mxwt_pconst),
      .din_2_rsci_biwt(din_2_rsci_biwt),
      .din_2_rsci_bdwt(din_2_rsci_bdwt)
    );
  assign din_2_rsci_douta_d_mxwt = din_2_rsci_douta_d_mxwt_pconst;
  assign din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_2_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1 (
  clk, rst, din_1_rsci_douta_d, din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_1_rsci_oswt, din_1_rsci_douta_d_mxwt, din_1_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_1_rsci_douta_d;
  output din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_1_rsci_oswt;
  output [15:0] din_1_rsci_douta_d_mxwt;
  input din_1_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_1_rsci_biwt;
  wire din_1_rsci_bdwt;
  wire [15:0] din_1_rsci_douta_d_mxwt_pconst;
  wire din_1_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1_din_1_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1_din_1_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_1_rsci_oswt(din_1_rsci_oswt),
      .din_1_rsci_biwt(din_1_rsci_biwt),
      .din_1_rsci_bdwt(din_1_rsci_bdwt),
      .din_1_rsci_biwt_pff(din_1_rsci_biwt_iff),
      .din_1_rsci_oswt_pff(din_1_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1_din_1_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1_din_1_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_1_rsci_douta_d(din_1_rsci_douta_d),
      .din_1_rsci_douta_d_mxwt(din_1_rsci_douta_d_mxwt_pconst),
      .din_1_rsci_biwt(din_1_rsci_biwt),
      .din_1_rsci_bdwt(din_1_rsci_bdwt)
    );
  assign din_1_rsci_douta_d_mxwt = din_1_rsci_douta_d_mxwt_pconst;
  assign din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_1_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1 (
  clk, rst, din_0_rsci_douta_d, din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      din_0_rsci_oswt, din_0_rsci_douta_d_mxwt, core_wten, din_0_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_0_rsci_douta_d;
  output din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input din_0_rsci_oswt;
  output [15:0] din_0_rsci_douta_d_mxwt;
  input core_wten;
  input din_0_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_0_rsci_biwt;
  wire din_0_rsci_bdwt;
  wire [15:0] din_0_rsci_douta_d_mxwt_pconst;
  wire din_0_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1_din_0_rsc_wait_ctrl READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1_din_0_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .din_0_rsci_oswt(din_0_rsci_oswt),
      .core_wten(core_wten),
      .din_0_rsci_biwt(din_0_rsci_biwt),
      .din_0_rsci_bdwt(din_0_rsci_bdwt),
      .din_0_rsci_biwt_pff(din_0_rsci_biwt_iff),
      .din_0_rsci_oswt_pff(din_0_rsci_oswt_pff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1_din_0_rsc_wait_dp READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1_din_0_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_0_rsci_douta_d(din_0_rsci_douta_d),
      .din_0_rsci_douta_d_mxwt(din_0_rsci_douta_d_mxwt_pconst),
      .din_0_rsci_biwt(din_0_rsci_biwt),
      .din_0_rsci_bdwt(din_0_rsci_bdwt)
    );
  assign din_0_rsci_douta_d_mxwt = din_0_rsci_douta_d_mxwt_pconst;
  assign din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_0_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj (
  clk, rst, dout_rsc_req_vz, core_wen, core_wten, dout_rsc_req_obj_oswt, dout_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_rsc_req_obj_oswt;
  output dout_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_rsc_req_obj_vd;
  wire dout_rsc_req_obj_biwt;
  wire dout_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_rsc_req_obj (
      .vd(dout_rsc_req_obj_vd),
      .vz(dout_rsc_req_vz)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
      WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj_dout_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsc_req_obj_oswt(dout_rsc_req_obj_oswt),
      .dout_rsc_req_obj_vd(dout_rsc_req_obj_vd),
      .dout_rsc_req_obj_biwt(dout_rsc_req_obj_biwt),
      .dout_rsc_req_obj_bdwt(dout_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj_dout_rsc_req_wait_dp WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj_dout_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_rsc_req_obj_oswt(dout_rsc_req_obj_oswt),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp),
      .dout_rsc_req_obj_biwt(dout_rsc_req_obj_biwt),
      .dout_rsc_req_obj_bdwt(dout_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_rls_obj (
  dout_rsc_rls_lz, core_wten, dout_rsc_rls_obj_iswt0
);
  output dout_rsc_rls_lz;
  input core_wten;
  input dout_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_rsc_rls_obj (
      .ld(dout_rsc_rls_obj_ld_core_sct),
      .lz(dout_rsc_rls_lz)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
      WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_rsc_rls_obj_iswt0(dout_rsc_rls_obj_iswt0),
      .dout_rsc_rls_obj_ld_core_sct(dout_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1 (
  dout_rsci_addra_d, dout_rsci_addrb_d, dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_rsci_addra_d_core, dout_rsci_addrb_d_core, dout_rsci_iswt0_pff, core_wten_pff
);
  output [6:0] dout_rsci_addra_d;
  output [6:0] dout_rsci_addrb_d;
  output dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input [6:0] dout_rsci_addra_d_core;
  input [6:0] dout_rsci_addrb_d_core;
  input dout_rsci_iswt0_pff;
  input core_wten_pff;


  // Interconnect Declarations
  wire dout_rsci_addra_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_dout_rsc_wait_ctrl WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_dout_rsc_wait_ctrl_inst
      (
      .dout_rsci_addra_d_core_sct_pff(dout_rsci_addra_d_core_sct_iff),
      .dout_rsci_iswt0_pff(dout_rsci_iswt0_pff),
      .core_wten_pff(core_wten_pff)
    );
  assign dout_rsci_addra_d = {(~ dout_rsci_addra_d_core_sct_iff) , (dout_rsci_addra_d_core[5:0])};
  assign dout_rsci_addrb_d = {(~ dout_rsci_addra_d_core_sct_iff) , (dout_rsci_addrb_d_core[5:0])};
  assign dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_rsci_addra_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, core_wen, din_rsci_oswt, din_rsci_wen_comp,
      din_rsci_d_mxwt, core_wten
);
  input clk;
  input rst;
  input [63:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  input core_wen;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [63:0] din_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire din_rsci_ld_core_sct;
  wire din_rsci_vd;
  wire [63:0] din_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_wait_v1 #(.rscid(32'sd95),
  .width(32'sd64)) din_rsci (
      .ld(din_rsci_ld_core_sct),
      .vd(din_rsci_vd),
      .d(din_rsci_d),
      .lz(din_rsc_lz),
      .vz(din_rsc_vz),
      .z(din_rsc_z)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci_din_wait_ctrl WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci_din_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .din_rsci_oswt(din_rsci_oswt),
      .core_wten(core_wten),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_ld_core_sct(din_rsci_ld_core_sct),
      .din_rsci_vd(din_rsci_vd)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci_din_wait_dp WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci_din_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_d_mxwt(din_rsci_d_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_d(din_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj (
  clk, rst, din_rsc_req_vz, core_wen, core_wten, din_rsc_req_obj_oswt, din_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_rsc_req_obj_oswt;
  output din_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_rsc_req_obj_vd;
  wire din_rsc_req_obj_biwt;
  wire din_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_rsc_req_obj (
      .vd(din_rsc_req_obj_vd),
      .vz(din_rsc_req_vz)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj_din_rsc_req_wait_ctrl
      READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj_din_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_rsc_req_obj_oswt(din_rsc_req_obj_oswt),
      .din_rsc_req_obj_vd(din_rsc_req_obj_vd),
      .din_rsc_req_obj_biwt(din_rsc_req_obj_biwt),
      .din_rsc_req_obj_bdwt(din_rsc_req_obj_bdwt)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj_din_rsc_req_wait_dp READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj_din_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_req_obj_oswt(din_rsc_req_obj_oswt),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp),
      .din_rsc_req_obj_biwt(din_rsc_req_obj_biwt),
      .din_rsc_req_obj_bdwt(din_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_rls_obj (
  din_rsc_rls_lz, core_wten, din_rsc_rls_obj_iswt0
);
  output din_rsc_rls_lz;
  input core_wten;
  input din_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_rsc_rls_obj (
      .ld(din_rsc_rls_obj_ld_core_sct),
      .lz(din_rsc_rls_lz)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
      READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_rls_obj_din_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_rsc_rls_obj_iswt0(din_rsc_rls_obj_iswt0),
      .din_rsc_rls_obj_ld_core_sct(din_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci (
  clk, rst, dout_rsc_z, dout_rsc_vz, dout_rsc_lz, core_wen, core_wten, dout_rsci_oswt,
      dout_rsci_wen_comp, dout_rsci_d
);
  input clk;
  input rst;
  output [63:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;
  input core_wen;
  input core_wten;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input [63:0] dout_rsci_d;


  // Interconnect Declarations
  wire dout_rsci_biwt;
  wire dout_rsci_bdwt;
  wire dout_rsci_ld_core_sct;
  wire dout_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  mgc_out_stdreg_wait_v1 #(.rscid(32'sd99),
  .width(32'sd64)) dout_rsci (
      .ld(dout_rsci_ld_core_sct),
      .vd(dout_rsci_vd),
      .d(dout_rsci_d),
      .lz(dout_rsc_lz),
      .vz(dout_rsc_vz),
      .z(dout_rsc_z)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci_dout_wait_ctrl READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci_dout_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_ld_core_sct(dout_rsci_ld_core_sct),
      .dout_rsci_vd(dout_rsci_vd)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci_dout_wait_dp READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci_dout_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1 (
  clk, rst, din_rsci_addra_d, din_rsci_addrb_d, din_rsci_douta_d, din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, din_rsci_oswt, din_rsci_addra_d_core, din_rsci_addrb_d_core, din_rsci_douta_d_mxwt,
      core_wten, din_rsci_oswt_pff
);
  input clk;
  input rst;
  output [6:0] din_rsci_addra_d;
  output [6:0] din_rsci_addrb_d;
  input [63:0] din_rsci_douta_d;
  output din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input din_rsci_oswt;
  input [6:0] din_rsci_addra_d_core;
  input [6:0] din_rsci_addrb_d_core;
  output [63:0] din_rsci_douta_d_mxwt;
  input core_wten;
  input din_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire [6:0] din_rsci_addra_d_reg;
  wire din_rsci_biwt_iff;
  wire [6:0] din_rsci_addrb_d_reg;


  // Interconnect Declarations for Component Instantiations 
  wire [6:0] nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addra_d_core;
  assign nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addra_d_core
      = {1'b0 , (din_rsci_addra_d_core[5:0])};
  wire [6:0] nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addrb_d_core;
  assign nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addrb_d_core
      = {1'b0 , (din_rsci_addrb_d_core[5:0])};
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_ctrl READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .din_rsci_oswt(din_rsci_oswt),
      .core_wten(core_wten),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_biwt_pff(din_rsci_biwt_iff),
      .din_rsci_oswt_pff(din_rsci_oswt_pff)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_dp READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsci_addra_d(din_rsci_addra_d_reg),
      .din_rsci_addrb_d(din_rsci_addrb_d_reg),
      .din_rsci_douta_d(din_rsci_douta_d),
      .din_rsci_addra_d_core(nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addra_d_core[6:0]),
      .din_rsci_addrb_d_core(nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addrb_d_core[6:0]),
      .din_rsci_douta_d_mxwt(din_rsci_douta_d_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_biwt_pff(din_rsci_biwt_iff)
    );
  assign din_rsci_addra_d = din_rsci_addra_d_reg;
  assign din_rsci_addrb_d = din_rsci_addrb_d_reg;
  assign din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core_output_rsci
// ------------------------------------------------------------------


module systolic_array_core_output_rsci (
  clk, rst, output_rsc_z, output_rsc_vz, output_rsc_lz, core_wen, core_wten, output_rsci_oswt,
      output_rsci_wen_comp, output_rsci_d
);
  input clk;
  input rst;
  output [1023:0] output_rsc_z;
  input output_rsc_vz;
  output output_rsc_lz;
  input core_wen;
  input core_wten;
  input output_rsci_oswt;
  output output_rsci_wen_comp;
  input [1023:0] output_rsci_d;


  // Interconnect Declarations
  wire output_rsci_biwt;
  wire output_rsci_bdwt;
  wire output_rsci_ld_core_sct;
  wire output_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  mgc_out_stdreg_wait_v1 #(.rscid(32'sd106),
  .width(32'sd1024)) output_rsci (
      .ld(output_rsci_ld_core_sct),
      .vd(output_rsci_vd),
      .d(output_rsci_d),
      .lz(output_rsc_lz),
      .vz(output_rsc_vz),
      .z(output_rsc_z)
    );
  systolic_array_core_output_rsci_output_wait_ctrl systolic_array_core_output_rsci_output_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .output_rsci_oswt(output_rsci_oswt),
      .output_rsci_biwt(output_rsci_biwt),
      .output_rsci_bdwt(output_rsci_bdwt),
      .output_rsci_ld_core_sct(output_rsci_ld_core_sct),
      .output_rsci_vd(output_rsci_vd)
    );
  systolic_array_core_output_rsci_output_wait_dp systolic_array_core_output_rsci_output_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .output_rsci_oswt(output_rsci_oswt),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .output_rsci_biwt(output_rsci_biwt),
      .output_rsci_bdwt(output_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core_weight_rsci
// ------------------------------------------------------------------


module systolic_array_core_weight_rsci (
  clk, rst, weight_rsc_z, weight_rsc_vz, weight_rsc_lz, core_wen, core_wten, weight_rsci_oswt,
      weight_rsci_wen_comp, weight_rsci_d_mxwt
);
  input clk;
  input rst;
  input [63:0] weight_rsc_z;
  input weight_rsc_vz;
  output weight_rsc_lz;
  input core_wen;
  input core_wten;
  input weight_rsci_oswt;
  output weight_rsci_wen_comp;
  output [31:0] weight_rsci_d_mxwt;


  // Interconnect Declarations
  wire weight_rsci_biwt;
  wire weight_rsci_bdwt;
  wire weight_rsci_ld_core_sct;
  wire weight_rsci_vd;
  wire [63:0] weight_rsci_d;
  wire [31:0] weight_rsci_d_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_wait_v1 #(.rscid(32'sd105),
  .width(32'sd64)) weight_rsci (
      .ld(weight_rsci_ld_core_sct),
      .vd(weight_rsci_vd),
      .d(weight_rsci_d),
      .lz(weight_rsc_lz),
      .vz(weight_rsc_vz),
      .z(weight_rsc_z)
    );
  systolic_array_core_weight_rsci_weight_wait_ctrl systolic_array_core_weight_rsci_weight_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .weight_rsci_oswt(weight_rsci_oswt),
      .weight_rsci_biwt(weight_rsci_biwt),
      .weight_rsci_bdwt(weight_rsci_bdwt),
      .weight_rsci_ld_core_sct(weight_rsci_ld_core_sct),
      .weight_rsci_vd(weight_rsci_vd)
    );
  systolic_array_core_weight_rsci_weight_wait_dp systolic_array_core_weight_rsci_weight_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .weight_rsci_oswt(weight_rsci_oswt),
      .weight_rsci_wen_comp(weight_rsci_wen_comp),
      .weight_rsci_d_mxwt(weight_rsci_d_mxwt_pconst),
      .weight_rsci_biwt(weight_rsci_biwt),
      .weight_rsci_bdwt(weight_rsci_bdwt),
      .weight_rsci_d(weight_rsci_d)
    );
  assign weight_rsci_d_mxwt = weight_rsci_d_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core_input_rsci
// ------------------------------------------------------------------


module systolic_array_core_input_rsci (
  clk, rst, input_rsc_z, input_rsc_vz, input_rsc_lz, core_wen, input_rsci_oswt, input_rsci_wen_comp,
      input_rsci_d_mxwt, core_wten
);
  input clk;
  input rst;
  input [511:0] input_rsc_z;
  input input_rsc_vz;
  output input_rsc_lz;
  input core_wen;
  input input_rsci_oswt;
  output input_rsci_wen_comp;
  output [255:0] input_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire input_rsci_biwt;
  wire input_rsci_bdwt;
  wire input_rsci_ld_core_sct;
  wire input_rsci_vd;
  wire [511:0] input_rsci_d;
  wire [255:0] input_rsci_d_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_wait_v1 #(.rscid(32'sd104),
  .width(32'sd512)) input_rsci (
      .ld(input_rsci_ld_core_sct),
      .vd(input_rsci_vd),
      .d(input_rsci_d),
      .lz(input_rsc_lz),
      .vz(input_rsc_vz),
      .z(input_rsc_z)
    );
  systolic_array_core_input_rsci_input_wait_ctrl systolic_array_core_input_rsci_input_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .input_rsci_oswt(input_rsci_oswt),
      .core_wten(core_wten),
      .input_rsci_biwt(input_rsci_biwt),
      .input_rsci_bdwt(input_rsci_bdwt),
      .input_rsci_ld_core_sct(input_rsci_ld_core_sct),
      .input_rsci_vd(input_rsci_vd)
    );
  systolic_array_core_input_rsci_input_wait_dp systolic_array_core_input_rsci_input_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_rsci_oswt(input_rsci_oswt),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .input_rsci_d_mxwt(input_rsci_d_mxwt_pconst),
      .input_rsci_biwt(input_rsci_biwt),
      .input_rsci_bdwt(input_rsci_bdwt),
      .input_rsci_d(input_rsci_d)
    );
  assign input_rsci_d_mxwt = input_rsci_d_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj (
  clk, rst, dout_0_rsc_req_vz, core_wen, core_wten, dout_0_rsc_req_obj_oswt, dout_0_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_0_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_0_rsc_req_obj_oswt;
  output dout_0_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_0_rsc_req_obj_vd;
  wire dout_0_rsc_req_obj_biwt;
  wire dout_0_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_0_rsc_req_obj (
      .vd(dout_0_rsc_req_obj_vd),
      .vz(dout_0_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_0_rsc_req_obj_oswt(dout_0_rsc_req_obj_oswt),
      .dout_0_rsc_req_obj_vd(dout_0_rsc_req_obj_vd),
      .dout_0_rsc_req_obj_biwt(dout_0_rsc_req_obj_biwt),
      .dout_0_rsc_req_obj_bdwt(dout_0_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj_dout_0_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_0_rsc_req_obj_oswt(dout_0_rsc_req_obj_oswt),
      .dout_0_rsc_req_obj_wen_comp(dout_0_rsc_req_obj_wen_comp),
      .dout_0_rsc_req_obj_biwt(dout_0_rsc_req_obj_biwt),
      .dout_0_rsc_req_obj_bdwt(dout_0_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj (
  clk, rst, dout_1_rsc_req_vz, core_wen, core_wten, dout_1_rsc_req_obj_oswt, dout_1_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_1_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_1_rsc_req_obj_oswt;
  output dout_1_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_1_rsc_req_obj_vd;
  wire dout_1_rsc_req_obj_biwt;
  wire dout_1_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_1_rsc_req_obj (
      .vd(dout_1_rsc_req_obj_vd),
      .vz(dout_1_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_1_rsc_req_obj_oswt(dout_1_rsc_req_obj_oswt),
      .dout_1_rsc_req_obj_vd(dout_1_rsc_req_obj_vd),
      .dout_1_rsc_req_obj_biwt(dout_1_rsc_req_obj_biwt),
      .dout_1_rsc_req_obj_bdwt(dout_1_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj_dout_1_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_1_rsc_req_obj_oswt(dout_1_rsc_req_obj_oswt),
      .dout_1_rsc_req_obj_wen_comp(dout_1_rsc_req_obj_wen_comp),
      .dout_1_rsc_req_obj_biwt(dout_1_rsc_req_obj_biwt),
      .dout_1_rsc_req_obj_bdwt(dout_1_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj (
  clk, rst, dout_2_rsc_req_vz, core_wen, core_wten, dout_2_rsc_req_obj_oswt, dout_2_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_2_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_2_rsc_req_obj_oswt;
  output dout_2_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_2_rsc_req_obj_vd;
  wire dout_2_rsc_req_obj_biwt;
  wire dout_2_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_2_rsc_req_obj (
      .vd(dout_2_rsc_req_obj_vd),
      .vz(dout_2_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_2_rsc_req_obj_oswt(dout_2_rsc_req_obj_oswt),
      .dout_2_rsc_req_obj_vd(dout_2_rsc_req_obj_vd),
      .dout_2_rsc_req_obj_biwt(dout_2_rsc_req_obj_biwt),
      .dout_2_rsc_req_obj_bdwt(dout_2_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj_dout_2_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_2_rsc_req_obj_oswt(dout_2_rsc_req_obj_oswt),
      .dout_2_rsc_req_obj_wen_comp(dout_2_rsc_req_obj_wen_comp),
      .dout_2_rsc_req_obj_biwt(dout_2_rsc_req_obj_biwt),
      .dout_2_rsc_req_obj_bdwt(dout_2_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj (
  clk, rst, dout_3_rsc_req_vz, core_wen, core_wten, dout_3_rsc_req_obj_oswt, dout_3_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_3_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_3_rsc_req_obj_oswt;
  output dout_3_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_3_rsc_req_obj_vd;
  wire dout_3_rsc_req_obj_biwt;
  wire dout_3_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_3_rsc_req_obj (
      .vd(dout_3_rsc_req_obj_vd),
      .vz(dout_3_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_3_rsc_req_obj_oswt(dout_3_rsc_req_obj_oswt),
      .dout_3_rsc_req_obj_vd(dout_3_rsc_req_obj_vd),
      .dout_3_rsc_req_obj_biwt(dout_3_rsc_req_obj_biwt),
      .dout_3_rsc_req_obj_bdwt(dout_3_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj_dout_3_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_3_rsc_req_obj_oswt(dout_3_rsc_req_obj_oswt),
      .dout_3_rsc_req_obj_wen_comp(dout_3_rsc_req_obj_wen_comp),
      .dout_3_rsc_req_obj_biwt(dout_3_rsc_req_obj_biwt),
      .dout_3_rsc_req_obj_bdwt(dout_3_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj (
  clk, rst, dout_4_rsc_req_vz, core_wen, core_wten, dout_4_rsc_req_obj_oswt, dout_4_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_4_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_4_rsc_req_obj_oswt;
  output dout_4_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_4_rsc_req_obj_vd;
  wire dout_4_rsc_req_obj_biwt;
  wire dout_4_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_4_rsc_req_obj (
      .vd(dout_4_rsc_req_obj_vd),
      .vz(dout_4_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_4_rsc_req_obj_oswt(dout_4_rsc_req_obj_oswt),
      .dout_4_rsc_req_obj_vd(dout_4_rsc_req_obj_vd),
      .dout_4_rsc_req_obj_biwt(dout_4_rsc_req_obj_biwt),
      .dout_4_rsc_req_obj_bdwt(dout_4_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj_dout_4_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_4_rsc_req_obj_oswt(dout_4_rsc_req_obj_oswt),
      .dout_4_rsc_req_obj_wen_comp(dout_4_rsc_req_obj_wen_comp),
      .dout_4_rsc_req_obj_biwt(dout_4_rsc_req_obj_biwt),
      .dout_4_rsc_req_obj_bdwt(dout_4_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj (
  clk, rst, dout_5_rsc_req_vz, core_wen, core_wten, dout_5_rsc_req_obj_oswt, dout_5_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_5_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_5_rsc_req_obj_oswt;
  output dout_5_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_5_rsc_req_obj_vd;
  wire dout_5_rsc_req_obj_biwt;
  wire dout_5_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_5_rsc_req_obj (
      .vd(dout_5_rsc_req_obj_vd),
      .vz(dout_5_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_5_rsc_req_obj_oswt(dout_5_rsc_req_obj_oswt),
      .dout_5_rsc_req_obj_vd(dout_5_rsc_req_obj_vd),
      .dout_5_rsc_req_obj_biwt(dout_5_rsc_req_obj_biwt),
      .dout_5_rsc_req_obj_bdwt(dout_5_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj_dout_5_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_5_rsc_req_obj_oswt(dout_5_rsc_req_obj_oswt),
      .dout_5_rsc_req_obj_wen_comp(dout_5_rsc_req_obj_wen_comp),
      .dout_5_rsc_req_obj_biwt(dout_5_rsc_req_obj_biwt),
      .dout_5_rsc_req_obj_bdwt(dout_5_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj (
  clk, rst, dout_6_rsc_req_vz, core_wen, core_wten, dout_6_rsc_req_obj_oswt, dout_6_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_6_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_6_rsc_req_obj_oswt;
  output dout_6_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_6_rsc_req_obj_vd;
  wire dout_6_rsc_req_obj_biwt;
  wire dout_6_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_6_rsc_req_obj (
      .vd(dout_6_rsc_req_obj_vd),
      .vz(dout_6_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_6_rsc_req_obj_oswt(dout_6_rsc_req_obj_oswt),
      .dout_6_rsc_req_obj_vd(dout_6_rsc_req_obj_vd),
      .dout_6_rsc_req_obj_biwt(dout_6_rsc_req_obj_biwt),
      .dout_6_rsc_req_obj_bdwt(dout_6_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj_dout_6_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_6_rsc_req_obj_oswt(dout_6_rsc_req_obj_oswt),
      .dout_6_rsc_req_obj_wen_comp(dout_6_rsc_req_obj_wen_comp),
      .dout_6_rsc_req_obj_biwt(dout_6_rsc_req_obj_biwt),
      .dout_6_rsc_req_obj_bdwt(dout_6_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj (
  clk, rst, dout_7_rsc_req_vz, core_wen, core_wten, dout_7_rsc_req_obj_oswt, dout_7_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_7_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_7_rsc_req_obj_oswt;
  output dout_7_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_7_rsc_req_obj_vd;
  wire dout_7_rsc_req_obj_biwt;
  wire dout_7_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_7_rsc_req_obj (
      .vd(dout_7_rsc_req_obj_vd),
      .vz(dout_7_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_7_rsc_req_obj_oswt(dout_7_rsc_req_obj_oswt),
      .dout_7_rsc_req_obj_vd(dout_7_rsc_req_obj_vd),
      .dout_7_rsc_req_obj_biwt(dout_7_rsc_req_obj_biwt),
      .dout_7_rsc_req_obj_bdwt(dout_7_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj_dout_7_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_7_rsc_req_obj_oswt(dout_7_rsc_req_obj_oswt),
      .dout_7_rsc_req_obj_wen_comp(dout_7_rsc_req_obj_wen_comp),
      .dout_7_rsc_req_obj_biwt(dout_7_rsc_req_obj_biwt),
      .dout_7_rsc_req_obj_bdwt(dout_7_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj (
  clk, rst, dout_8_rsc_req_vz, core_wen, core_wten, dout_8_rsc_req_obj_oswt, dout_8_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_8_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_8_rsc_req_obj_oswt;
  output dout_8_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_8_rsc_req_obj_vd;
  wire dout_8_rsc_req_obj_biwt;
  wire dout_8_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_8_rsc_req_obj (
      .vd(dout_8_rsc_req_obj_vd),
      .vz(dout_8_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_8_rsc_req_obj_oswt(dout_8_rsc_req_obj_oswt),
      .dout_8_rsc_req_obj_vd(dout_8_rsc_req_obj_vd),
      .dout_8_rsc_req_obj_biwt(dout_8_rsc_req_obj_biwt),
      .dout_8_rsc_req_obj_bdwt(dout_8_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj_dout_8_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_8_rsc_req_obj_oswt(dout_8_rsc_req_obj_oswt),
      .dout_8_rsc_req_obj_wen_comp(dout_8_rsc_req_obj_wen_comp),
      .dout_8_rsc_req_obj_biwt(dout_8_rsc_req_obj_biwt),
      .dout_8_rsc_req_obj_bdwt(dout_8_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj (
  clk, rst, dout_9_rsc_req_vz, core_wen, core_wten, dout_9_rsc_req_obj_oswt, dout_9_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_9_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_9_rsc_req_obj_oswt;
  output dout_9_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_9_rsc_req_obj_vd;
  wire dout_9_rsc_req_obj_biwt;
  wire dout_9_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_9_rsc_req_obj (
      .vd(dout_9_rsc_req_obj_vd),
      .vz(dout_9_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_9_rsc_req_obj_oswt(dout_9_rsc_req_obj_oswt),
      .dout_9_rsc_req_obj_vd(dout_9_rsc_req_obj_vd),
      .dout_9_rsc_req_obj_biwt(dout_9_rsc_req_obj_biwt),
      .dout_9_rsc_req_obj_bdwt(dout_9_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj_dout_9_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_9_rsc_req_obj_oswt(dout_9_rsc_req_obj_oswt),
      .dout_9_rsc_req_obj_wen_comp(dout_9_rsc_req_obj_wen_comp),
      .dout_9_rsc_req_obj_biwt(dout_9_rsc_req_obj_biwt),
      .dout_9_rsc_req_obj_bdwt(dout_9_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj (
  clk, rst, dout_10_rsc_req_vz, core_wen, core_wten, dout_10_rsc_req_obj_oswt, dout_10_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_10_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_10_rsc_req_obj_oswt;
  output dout_10_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_10_rsc_req_obj_vd;
  wire dout_10_rsc_req_obj_biwt;
  wire dout_10_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_10_rsc_req_obj (
      .vd(dout_10_rsc_req_obj_vd),
      .vz(dout_10_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_10_rsc_req_obj_oswt(dout_10_rsc_req_obj_oswt),
      .dout_10_rsc_req_obj_vd(dout_10_rsc_req_obj_vd),
      .dout_10_rsc_req_obj_biwt(dout_10_rsc_req_obj_biwt),
      .dout_10_rsc_req_obj_bdwt(dout_10_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj_dout_10_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_10_rsc_req_obj_oswt(dout_10_rsc_req_obj_oswt),
      .dout_10_rsc_req_obj_wen_comp(dout_10_rsc_req_obj_wen_comp),
      .dout_10_rsc_req_obj_biwt(dout_10_rsc_req_obj_biwt),
      .dout_10_rsc_req_obj_bdwt(dout_10_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj (
  clk, rst, dout_11_rsc_req_vz, core_wen, core_wten, dout_11_rsc_req_obj_oswt, dout_11_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_11_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_11_rsc_req_obj_oswt;
  output dout_11_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_11_rsc_req_obj_vd;
  wire dout_11_rsc_req_obj_biwt;
  wire dout_11_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_11_rsc_req_obj (
      .vd(dout_11_rsc_req_obj_vd),
      .vz(dout_11_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_11_rsc_req_obj_oswt(dout_11_rsc_req_obj_oswt),
      .dout_11_rsc_req_obj_vd(dout_11_rsc_req_obj_vd),
      .dout_11_rsc_req_obj_biwt(dout_11_rsc_req_obj_biwt),
      .dout_11_rsc_req_obj_bdwt(dout_11_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj_dout_11_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_11_rsc_req_obj_oswt(dout_11_rsc_req_obj_oswt),
      .dout_11_rsc_req_obj_wen_comp(dout_11_rsc_req_obj_wen_comp),
      .dout_11_rsc_req_obj_biwt(dout_11_rsc_req_obj_biwt),
      .dout_11_rsc_req_obj_bdwt(dout_11_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj (
  clk, rst, dout_12_rsc_req_vz, core_wen, core_wten, dout_12_rsc_req_obj_oswt, dout_12_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_12_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_12_rsc_req_obj_oswt;
  output dout_12_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_12_rsc_req_obj_vd;
  wire dout_12_rsc_req_obj_biwt;
  wire dout_12_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_12_rsc_req_obj (
      .vd(dout_12_rsc_req_obj_vd),
      .vz(dout_12_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_12_rsc_req_obj_oswt(dout_12_rsc_req_obj_oswt),
      .dout_12_rsc_req_obj_vd(dout_12_rsc_req_obj_vd),
      .dout_12_rsc_req_obj_biwt(dout_12_rsc_req_obj_biwt),
      .dout_12_rsc_req_obj_bdwt(dout_12_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj_dout_12_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_12_rsc_req_obj_oswt(dout_12_rsc_req_obj_oswt),
      .dout_12_rsc_req_obj_wen_comp(dout_12_rsc_req_obj_wen_comp),
      .dout_12_rsc_req_obj_biwt(dout_12_rsc_req_obj_biwt),
      .dout_12_rsc_req_obj_bdwt(dout_12_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj (
  clk, rst, dout_13_rsc_req_vz, core_wen, core_wten, dout_13_rsc_req_obj_oswt, dout_13_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_13_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_13_rsc_req_obj_oswt;
  output dout_13_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_13_rsc_req_obj_vd;
  wire dout_13_rsc_req_obj_biwt;
  wire dout_13_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_13_rsc_req_obj (
      .vd(dout_13_rsc_req_obj_vd),
      .vz(dout_13_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_13_rsc_req_obj_oswt(dout_13_rsc_req_obj_oswt),
      .dout_13_rsc_req_obj_vd(dout_13_rsc_req_obj_vd),
      .dout_13_rsc_req_obj_biwt(dout_13_rsc_req_obj_biwt),
      .dout_13_rsc_req_obj_bdwt(dout_13_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj_dout_13_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_13_rsc_req_obj_oswt(dout_13_rsc_req_obj_oswt),
      .dout_13_rsc_req_obj_wen_comp(dout_13_rsc_req_obj_wen_comp),
      .dout_13_rsc_req_obj_biwt(dout_13_rsc_req_obj_biwt),
      .dout_13_rsc_req_obj_bdwt(dout_13_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj (
  clk, rst, dout_14_rsc_req_vz, core_wen, core_wten, dout_14_rsc_req_obj_oswt, dout_14_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_14_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_14_rsc_req_obj_oswt;
  output dout_14_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_14_rsc_req_obj_vd;
  wire dout_14_rsc_req_obj_biwt;
  wire dout_14_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_14_rsc_req_obj (
      .vd(dout_14_rsc_req_obj_vd),
      .vz(dout_14_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_14_rsc_req_obj_oswt(dout_14_rsc_req_obj_oswt),
      .dout_14_rsc_req_obj_vd(dout_14_rsc_req_obj_vd),
      .dout_14_rsc_req_obj_biwt(dout_14_rsc_req_obj_biwt),
      .dout_14_rsc_req_obj_bdwt(dout_14_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj_dout_14_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_14_rsc_req_obj_oswt(dout_14_rsc_req_obj_oswt),
      .dout_14_rsc_req_obj_wen_comp(dout_14_rsc_req_obj_wen_comp),
      .dout_14_rsc_req_obj_biwt(dout_14_rsc_req_obj_biwt),
      .dout_14_rsc_req_obj_bdwt(dout_14_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj (
  clk, rst, dout_15_rsc_req_vz, core_wen, core_wten, dout_15_rsc_req_obj_oswt, dout_15_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input dout_15_rsc_req_vz;
  input core_wen;
  input core_wten;
  input dout_15_rsc_req_obj_oswt;
  output dout_15_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_15_rsc_req_obj_vd;
  wire dout_15_rsc_req_obj_biwt;
  wire dout_15_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) dout_15_rsc_req_obj (
      .vd(dout_15_rsc_req_obj_vd),
      .vz(dout_15_rsc_req_vz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_15_rsc_req_obj_oswt(dout_15_rsc_req_obj_oswt),
      .dout_15_rsc_req_obj_vd(dout_15_rsc_req_obj_vd),
      .dout_15_rsc_req_obj_biwt(dout_15_rsc_req_obj_biwt),
      .dout_15_rsc_req_obj_bdwt(dout_15_rsc_req_obj_bdwt)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_dp
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj_dout_15_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_15_rsc_req_obj_oswt(dout_15_rsc_req_obj_oswt),
      .dout_15_rsc_req_obj_wen_comp(dout_15_rsc_req_obj_wen_comp),
      .dout_15_rsc_req_obj_biwt(dout_15_rsc_req_obj_biwt),
      .dout_15_rsc_req_obj_bdwt(dout_15_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_rls_obj (
  dout_0_rsc_rls_lz, core_wten, dout_0_rsc_rls_obj_iswt0
);
  output dout_0_rsc_rls_lz;
  input core_wten;
  input dout_0_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_0_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_0_rsc_rls_obj (
      .ld(dout_0_rsc_rls_obj_ld_core_sct),
      .lz(dout_0_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_rls_obj_dout_0_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_rls_obj_dout_0_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_0_rsc_rls_obj_iswt0(dout_0_rsc_rls_obj_iswt0),
      .dout_0_rsc_rls_obj_ld_core_sct(dout_0_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_rls_obj (
  dout_1_rsc_rls_lz, core_wten, dout_1_rsc_rls_obj_iswt0
);
  output dout_1_rsc_rls_lz;
  input core_wten;
  input dout_1_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_1_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_1_rsc_rls_obj (
      .ld(dout_1_rsc_rls_obj_ld_core_sct),
      .lz(dout_1_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_rls_obj_dout_1_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_rls_obj_dout_1_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_1_rsc_rls_obj_iswt0(dout_1_rsc_rls_obj_iswt0),
      .dout_1_rsc_rls_obj_ld_core_sct(dout_1_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_rls_obj (
  dout_2_rsc_rls_lz, core_wten, dout_2_rsc_rls_obj_iswt0
);
  output dout_2_rsc_rls_lz;
  input core_wten;
  input dout_2_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_2_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_2_rsc_rls_obj (
      .ld(dout_2_rsc_rls_obj_ld_core_sct),
      .lz(dout_2_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_rls_obj_dout_2_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_rls_obj_dout_2_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_2_rsc_rls_obj_iswt0(dout_2_rsc_rls_obj_iswt0),
      .dout_2_rsc_rls_obj_ld_core_sct(dout_2_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_rls_obj (
  dout_3_rsc_rls_lz, core_wten, dout_3_rsc_rls_obj_iswt0
);
  output dout_3_rsc_rls_lz;
  input core_wten;
  input dout_3_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_3_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_3_rsc_rls_obj (
      .ld(dout_3_rsc_rls_obj_ld_core_sct),
      .lz(dout_3_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_rls_obj_dout_3_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_rls_obj_dout_3_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_3_rsc_rls_obj_iswt0(dout_3_rsc_rls_obj_iswt0),
      .dout_3_rsc_rls_obj_ld_core_sct(dout_3_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_rls_obj (
  dout_4_rsc_rls_lz, core_wten, dout_4_rsc_rls_obj_iswt0
);
  output dout_4_rsc_rls_lz;
  input core_wten;
  input dout_4_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_4_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_4_rsc_rls_obj (
      .ld(dout_4_rsc_rls_obj_ld_core_sct),
      .lz(dout_4_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_rls_obj_dout_4_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_rls_obj_dout_4_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_4_rsc_rls_obj_iswt0(dout_4_rsc_rls_obj_iswt0),
      .dout_4_rsc_rls_obj_ld_core_sct(dout_4_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_rls_obj (
  dout_5_rsc_rls_lz, core_wten, dout_5_rsc_rls_obj_iswt0
);
  output dout_5_rsc_rls_lz;
  input core_wten;
  input dout_5_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_5_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_5_rsc_rls_obj (
      .ld(dout_5_rsc_rls_obj_ld_core_sct),
      .lz(dout_5_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_rls_obj_dout_5_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_rls_obj_dout_5_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_5_rsc_rls_obj_iswt0(dout_5_rsc_rls_obj_iswt0),
      .dout_5_rsc_rls_obj_ld_core_sct(dout_5_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_rls_obj (
  dout_6_rsc_rls_lz, core_wten, dout_6_rsc_rls_obj_iswt0
);
  output dout_6_rsc_rls_lz;
  input core_wten;
  input dout_6_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_6_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_6_rsc_rls_obj (
      .ld(dout_6_rsc_rls_obj_ld_core_sct),
      .lz(dout_6_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_rls_obj_dout_6_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_rls_obj_dout_6_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_6_rsc_rls_obj_iswt0(dout_6_rsc_rls_obj_iswt0),
      .dout_6_rsc_rls_obj_ld_core_sct(dout_6_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_rls_obj (
  dout_7_rsc_rls_lz, core_wten, dout_7_rsc_rls_obj_iswt0
);
  output dout_7_rsc_rls_lz;
  input core_wten;
  input dout_7_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_7_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_7_rsc_rls_obj (
      .ld(dout_7_rsc_rls_obj_ld_core_sct),
      .lz(dout_7_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_rls_obj_dout_7_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_rls_obj_dout_7_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_7_rsc_rls_obj_iswt0(dout_7_rsc_rls_obj_iswt0),
      .dout_7_rsc_rls_obj_ld_core_sct(dout_7_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_rls_obj (
  dout_8_rsc_rls_lz, core_wten, dout_8_rsc_rls_obj_iswt0
);
  output dout_8_rsc_rls_lz;
  input core_wten;
  input dout_8_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_8_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_8_rsc_rls_obj (
      .ld(dout_8_rsc_rls_obj_ld_core_sct),
      .lz(dout_8_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_rls_obj_dout_8_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_rls_obj_dout_8_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_8_rsc_rls_obj_iswt0(dout_8_rsc_rls_obj_iswt0),
      .dout_8_rsc_rls_obj_ld_core_sct(dout_8_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_rls_obj (
  dout_9_rsc_rls_lz, core_wten, dout_9_rsc_rls_obj_iswt0
);
  output dout_9_rsc_rls_lz;
  input core_wten;
  input dout_9_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_9_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_9_rsc_rls_obj (
      .ld(dout_9_rsc_rls_obj_ld_core_sct),
      .lz(dout_9_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_rls_obj_dout_9_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_rls_obj_dout_9_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_9_rsc_rls_obj_iswt0(dout_9_rsc_rls_obj_iswt0),
      .dout_9_rsc_rls_obj_ld_core_sct(dout_9_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_rls_obj (
  dout_10_rsc_rls_lz, core_wten, dout_10_rsc_rls_obj_iswt0
);
  output dout_10_rsc_rls_lz;
  input core_wten;
  input dout_10_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_10_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_10_rsc_rls_obj (
      .ld(dout_10_rsc_rls_obj_ld_core_sct),
      .lz(dout_10_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_rls_obj_dout_10_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_rls_obj_dout_10_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_10_rsc_rls_obj_iswt0(dout_10_rsc_rls_obj_iswt0),
      .dout_10_rsc_rls_obj_ld_core_sct(dout_10_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_rls_obj (
  dout_11_rsc_rls_lz, core_wten, dout_11_rsc_rls_obj_iswt0
);
  output dout_11_rsc_rls_lz;
  input core_wten;
  input dout_11_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_11_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_11_rsc_rls_obj (
      .ld(dout_11_rsc_rls_obj_ld_core_sct),
      .lz(dout_11_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_rls_obj_dout_11_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_rls_obj_dout_11_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_11_rsc_rls_obj_iswt0(dout_11_rsc_rls_obj_iswt0),
      .dout_11_rsc_rls_obj_ld_core_sct(dout_11_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_rls_obj (
  dout_12_rsc_rls_lz, core_wten, dout_12_rsc_rls_obj_iswt0
);
  output dout_12_rsc_rls_lz;
  input core_wten;
  input dout_12_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_12_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_12_rsc_rls_obj (
      .ld(dout_12_rsc_rls_obj_ld_core_sct),
      .lz(dout_12_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_rls_obj_dout_12_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_rls_obj_dout_12_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_12_rsc_rls_obj_iswt0(dout_12_rsc_rls_obj_iswt0),
      .dout_12_rsc_rls_obj_ld_core_sct(dout_12_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_rls_obj (
  dout_13_rsc_rls_lz, core_wten, dout_13_rsc_rls_obj_iswt0
);
  output dout_13_rsc_rls_lz;
  input core_wten;
  input dout_13_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_13_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_13_rsc_rls_obj (
      .ld(dout_13_rsc_rls_obj_ld_core_sct),
      .lz(dout_13_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_rls_obj_dout_13_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_rls_obj_dout_13_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_13_rsc_rls_obj_iswt0(dout_13_rsc_rls_obj_iswt0),
      .dout_13_rsc_rls_obj_ld_core_sct(dout_13_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_rls_obj (
  dout_14_rsc_rls_lz, core_wten, dout_14_rsc_rls_obj_iswt0
);
  output dout_14_rsc_rls_lz;
  input core_wten;
  input dout_14_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_14_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_14_rsc_rls_obj (
      .ld(dout_14_rsc_rls_obj_ld_core_sct),
      .lz(dout_14_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_rls_obj_dout_14_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_rls_obj_dout_14_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_14_rsc_rls_obj_iswt0(dout_14_rsc_rls_obj_iswt0),
      .dout_14_rsc_rls_obj_ld_core_sct(dout_14_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_rls_obj
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_rls_obj (
  dout_15_rsc_rls_lz, core_wten, dout_15_rsc_rls_obj_iswt0
);
  output dout_15_rsc_rls_lz;
  input core_wten;
  input dout_15_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_15_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) dout_15_rsc_rls_obj (
      .ld(dout_15_rsc_rls_obj_ld_core_sct),
      .lz(dout_15_rsc_rls_lz)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_rls_obj_dout_15_rsc_rls_wait_ctrl
      WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_rls_obj_dout_15_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_15_rsc_rls_obj_iswt0(dout_15_rsc_rls_obj_iswt0),
      .dout_15_rsc_rls_obj_ld_core_sct(dout_15_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1 (
  dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_15_rsci_iswt0
);
  output dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_15_rsci_iswt0;


  // Interconnect Declarations
  wire dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_dout_15_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_dout_15_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_15_rsci_iswt0(dout_15_rsci_iswt0),
      .dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1 (
  dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_14_rsci_iswt0
);
  output dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_14_rsci_iswt0;


  // Interconnect Declarations
  wire dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_dout_14_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_dout_14_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_14_rsci_iswt0(dout_14_rsci_iswt0),
      .dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1 (
  dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_13_rsci_iswt0
);
  output dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_13_rsci_iswt0;


  // Interconnect Declarations
  wire dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_dout_13_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_dout_13_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_13_rsci_iswt0(dout_13_rsci_iswt0),
      .dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1 (
  dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_12_rsci_iswt0
);
  output dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_12_rsci_iswt0;


  // Interconnect Declarations
  wire dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_dout_12_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_dout_12_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_12_rsci_iswt0(dout_12_rsci_iswt0),
      .dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1 (
  dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_11_rsci_iswt0
);
  output dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_11_rsci_iswt0;


  // Interconnect Declarations
  wire dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_dout_11_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_dout_11_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_11_rsci_iswt0(dout_11_rsci_iswt0),
      .dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1 (
  dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_10_rsci_iswt0
);
  output dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_10_rsci_iswt0;


  // Interconnect Declarations
  wire dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_dout_10_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_dout_10_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_10_rsci_iswt0(dout_10_rsci_iswt0),
      .dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1 (
  dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_9_rsci_iswt0
);
  output dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_9_rsci_iswt0;


  // Interconnect Declarations
  wire dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_dout_9_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_dout_9_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_9_rsci_iswt0(dout_9_rsci_iswt0),
      .dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1 (
  dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_8_rsci_iswt0
);
  output dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_8_rsci_iswt0;


  // Interconnect Declarations
  wire dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_dout_8_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_dout_8_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_8_rsci_iswt0(dout_8_rsci_iswt0),
      .dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1 (
  dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_7_rsci_iswt0
);
  output dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_7_rsci_iswt0;


  // Interconnect Declarations
  wire dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_dout_7_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_dout_7_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_7_rsci_iswt0(dout_7_rsci_iswt0),
      .dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1 (
  dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_6_rsci_iswt0
);
  output dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_6_rsci_iswt0;


  // Interconnect Declarations
  wire dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_dout_6_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_dout_6_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_6_rsci_iswt0(dout_6_rsci_iswt0),
      .dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1 (
  dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_5_rsci_iswt0
);
  output dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_5_rsci_iswt0;


  // Interconnect Declarations
  wire dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_dout_5_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_dout_5_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_5_rsci_iswt0(dout_5_rsci_iswt0),
      .dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1 (
  dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_4_rsci_iswt0
);
  output dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_4_rsci_iswt0;


  // Interconnect Declarations
  wire dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_dout_4_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_dout_4_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_4_rsci_iswt0(dout_4_rsci_iswt0),
      .dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1 (
  dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_3_rsci_iswt0
);
  output dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_3_rsci_iswt0;


  // Interconnect Declarations
  wire dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_dout_3_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_dout_3_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_3_rsci_iswt0(dout_3_rsci_iswt0),
      .dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1 (
  dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_2_rsci_iswt0
);
  output dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_2_rsci_iswt0;


  // Interconnect Declarations
  wire dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_dout_2_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_dout_2_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_2_rsci_iswt0(dout_2_rsci_iswt0),
      .dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1 (
  dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_1_rsci_iswt0
);
  output dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_1_rsci_iswt0;


  // Interconnect Declarations
  wire dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_dout_1_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_dout_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_1_rsci_iswt0(dout_1_rsci_iswt0),
      .dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1 (
  dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, core_wten, dout_0_rsci_iswt0
);
  output dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  input core_wten;
  input dout_0_rsci_iswt0;


  // Interconnect Declarations
  wire dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_dout_0_rsc_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_dout_0_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .dout_0_rsci_iswt0(dout_0_rsci_iswt0),
      .dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct(dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct)
    );
  assign dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, core_wen, din_rsci_oswt, din_rsci_wen_comp,
      din_rsci_d_mxwt, core_wten
);
  input clk;
  input rst;
  input [1023:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  input core_wen;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [1023:0] din_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire din_rsci_ld_core_sct;
  wire din_rsci_vd;
  wire [1023:0] din_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_wait_v1 #(.rscid(32'sd112),
  .width(32'sd1024)) din_rsci (
      .ld(din_rsci_ld_core_sct),
      .vd(din_rsci_vd),
      .d(din_rsci_d),
      .lz(din_rsc_lz),
      .vz(din_rsc_vz),
      .z(din_rsc_z)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci_din_wait_ctrl WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci_din_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .din_rsci_oswt(din_rsci_oswt),
      .core_wten(core_wten),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_ld_core_sct(din_rsci_ld_core_sct),
      .din_rsci_vd(din_rsci_vd)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci_din_wait_dp WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci_din_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_d_mxwt(din_rsci_d_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_d(din_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj (
  clk, rst, din_0_rsc_req_vz, core_wen, core_wten, din_0_rsc_req_obj_oswt, din_0_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_0_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_0_rsc_req_obj_oswt;
  output din_0_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_0_rsc_req_obj_vd;
  wire din_0_rsc_req_obj_biwt;
  wire din_0_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_0_rsc_req_obj (
      .vd(din_0_rsc_req_obj_vd),
      .vz(din_0_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj_din_0_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj_din_0_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_0_rsc_req_obj_oswt(din_0_rsc_req_obj_oswt),
      .din_0_rsc_req_obj_vd(din_0_rsc_req_obj_vd),
      .din_0_rsc_req_obj_biwt(din_0_rsc_req_obj_biwt),
      .din_0_rsc_req_obj_bdwt(din_0_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj_din_0_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj_din_0_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_0_rsc_req_obj_oswt(din_0_rsc_req_obj_oswt),
      .din_0_rsc_req_obj_wen_comp(din_0_rsc_req_obj_wen_comp),
      .din_0_rsc_req_obj_biwt(din_0_rsc_req_obj_biwt),
      .din_0_rsc_req_obj_bdwt(din_0_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj (
  clk, rst, din_1_rsc_req_vz, core_wen, core_wten, din_1_rsc_req_obj_oswt, din_1_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_1_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_1_rsc_req_obj_oswt;
  output din_1_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_1_rsc_req_obj_vd;
  wire din_1_rsc_req_obj_biwt;
  wire din_1_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_1_rsc_req_obj (
      .vd(din_1_rsc_req_obj_vd),
      .vz(din_1_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj_din_1_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj_din_1_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_1_rsc_req_obj_oswt(din_1_rsc_req_obj_oswt),
      .din_1_rsc_req_obj_vd(din_1_rsc_req_obj_vd),
      .din_1_rsc_req_obj_biwt(din_1_rsc_req_obj_biwt),
      .din_1_rsc_req_obj_bdwt(din_1_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj_din_1_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj_din_1_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_1_rsc_req_obj_oswt(din_1_rsc_req_obj_oswt),
      .din_1_rsc_req_obj_wen_comp(din_1_rsc_req_obj_wen_comp),
      .din_1_rsc_req_obj_biwt(din_1_rsc_req_obj_biwt),
      .din_1_rsc_req_obj_bdwt(din_1_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj (
  clk, rst, din_2_rsc_req_vz, core_wen, core_wten, din_2_rsc_req_obj_oswt, din_2_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_2_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_2_rsc_req_obj_oswt;
  output din_2_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_2_rsc_req_obj_vd;
  wire din_2_rsc_req_obj_biwt;
  wire din_2_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_2_rsc_req_obj (
      .vd(din_2_rsc_req_obj_vd),
      .vz(din_2_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj_din_2_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj_din_2_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_2_rsc_req_obj_oswt(din_2_rsc_req_obj_oswt),
      .din_2_rsc_req_obj_vd(din_2_rsc_req_obj_vd),
      .din_2_rsc_req_obj_biwt(din_2_rsc_req_obj_biwt),
      .din_2_rsc_req_obj_bdwt(din_2_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj_din_2_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj_din_2_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_2_rsc_req_obj_oswt(din_2_rsc_req_obj_oswt),
      .din_2_rsc_req_obj_wen_comp(din_2_rsc_req_obj_wen_comp),
      .din_2_rsc_req_obj_biwt(din_2_rsc_req_obj_biwt),
      .din_2_rsc_req_obj_bdwt(din_2_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj (
  clk, rst, din_3_rsc_req_vz, core_wen, core_wten, din_3_rsc_req_obj_oswt, din_3_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_3_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_3_rsc_req_obj_oswt;
  output din_3_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_3_rsc_req_obj_vd;
  wire din_3_rsc_req_obj_biwt;
  wire din_3_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_3_rsc_req_obj (
      .vd(din_3_rsc_req_obj_vd),
      .vz(din_3_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj_din_3_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj_din_3_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_3_rsc_req_obj_oswt(din_3_rsc_req_obj_oswt),
      .din_3_rsc_req_obj_vd(din_3_rsc_req_obj_vd),
      .din_3_rsc_req_obj_biwt(din_3_rsc_req_obj_biwt),
      .din_3_rsc_req_obj_bdwt(din_3_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj_din_3_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj_din_3_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_3_rsc_req_obj_oswt(din_3_rsc_req_obj_oswt),
      .din_3_rsc_req_obj_wen_comp(din_3_rsc_req_obj_wen_comp),
      .din_3_rsc_req_obj_biwt(din_3_rsc_req_obj_biwt),
      .din_3_rsc_req_obj_bdwt(din_3_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj (
  clk, rst, din_4_rsc_req_vz, core_wen, core_wten, din_4_rsc_req_obj_oswt, din_4_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_4_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_4_rsc_req_obj_oswt;
  output din_4_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_4_rsc_req_obj_vd;
  wire din_4_rsc_req_obj_biwt;
  wire din_4_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_4_rsc_req_obj (
      .vd(din_4_rsc_req_obj_vd),
      .vz(din_4_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj_din_4_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj_din_4_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_4_rsc_req_obj_oswt(din_4_rsc_req_obj_oswt),
      .din_4_rsc_req_obj_vd(din_4_rsc_req_obj_vd),
      .din_4_rsc_req_obj_biwt(din_4_rsc_req_obj_biwt),
      .din_4_rsc_req_obj_bdwt(din_4_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj_din_4_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj_din_4_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_4_rsc_req_obj_oswt(din_4_rsc_req_obj_oswt),
      .din_4_rsc_req_obj_wen_comp(din_4_rsc_req_obj_wen_comp),
      .din_4_rsc_req_obj_biwt(din_4_rsc_req_obj_biwt),
      .din_4_rsc_req_obj_bdwt(din_4_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj (
  clk, rst, din_5_rsc_req_vz, core_wen, core_wten, din_5_rsc_req_obj_oswt, din_5_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_5_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_5_rsc_req_obj_oswt;
  output din_5_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_5_rsc_req_obj_vd;
  wire din_5_rsc_req_obj_biwt;
  wire din_5_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_5_rsc_req_obj (
      .vd(din_5_rsc_req_obj_vd),
      .vz(din_5_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj_din_5_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj_din_5_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_5_rsc_req_obj_oswt(din_5_rsc_req_obj_oswt),
      .din_5_rsc_req_obj_vd(din_5_rsc_req_obj_vd),
      .din_5_rsc_req_obj_biwt(din_5_rsc_req_obj_biwt),
      .din_5_rsc_req_obj_bdwt(din_5_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj_din_5_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj_din_5_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_5_rsc_req_obj_oswt(din_5_rsc_req_obj_oswt),
      .din_5_rsc_req_obj_wen_comp(din_5_rsc_req_obj_wen_comp),
      .din_5_rsc_req_obj_biwt(din_5_rsc_req_obj_biwt),
      .din_5_rsc_req_obj_bdwt(din_5_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj (
  clk, rst, din_6_rsc_req_vz, core_wen, core_wten, din_6_rsc_req_obj_oswt, din_6_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_6_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_6_rsc_req_obj_oswt;
  output din_6_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_6_rsc_req_obj_vd;
  wire din_6_rsc_req_obj_biwt;
  wire din_6_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_6_rsc_req_obj (
      .vd(din_6_rsc_req_obj_vd),
      .vz(din_6_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj_din_6_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj_din_6_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_6_rsc_req_obj_oswt(din_6_rsc_req_obj_oswt),
      .din_6_rsc_req_obj_vd(din_6_rsc_req_obj_vd),
      .din_6_rsc_req_obj_biwt(din_6_rsc_req_obj_biwt),
      .din_6_rsc_req_obj_bdwt(din_6_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj_din_6_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj_din_6_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_6_rsc_req_obj_oswt(din_6_rsc_req_obj_oswt),
      .din_6_rsc_req_obj_wen_comp(din_6_rsc_req_obj_wen_comp),
      .din_6_rsc_req_obj_biwt(din_6_rsc_req_obj_biwt),
      .din_6_rsc_req_obj_bdwt(din_6_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj (
  clk, rst, din_7_rsc_req_vz, core_wen, core_wten, din_7_rsc_req_obj_oswt, din_7_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_7_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_7_rsc_req_obj_oswt;
  output din_7_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_7_rsc_req_obj_vd;
  wire din_7_rsc_req_obj_biwt;
  wire din_7_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_7_rsc_req_obj (
      .vd(din_7_rsc_req_obj_vd),
      .vz(din_7_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj_din_7_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj_din_7_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_7_rsc_req_obj_oswt(din_7_rsc_req_obj_oswt),
      .din_7_rsc_req_obj_vd(din_7_rsc_req_obj_vd),
      .din_7_rsc_req_obj_biwt(din_7_rsc_req_obj_biwt),
      .din_7_rsc_req_obj_bdwt(din_7_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj_din_7_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj_din_7_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_7_rsc_req_obj_oswt(din_7_rsc_req_obj_oswt),
      .din_7_rsc_req_obj_wen_comp(din_7_rsc_req_obj_wen_comp),
      .din_7_rsc_req_obj_biwt(din_7_rsc_req_obj_biwt),
      .din_7_rsc_req_obj_bdwt(din_7_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj (
  clk, rst, din_8_rsc_req_vz, core_wen, core_wten, din_8_rsc_req_obj_oswt, din_8_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_8_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_8_rsc_req_obj_oswt;
  output din_8_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_8_rsc_req_obj_vd;
  wire din_8_rsc_req_obj_biwt;
  wire din_8_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_8_rsc_req_obj (
      .vd(din_8_rsc_req_obj_vd),
      .vz(din_8_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj_din_8_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj_din_8_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_8_rsc_req_obj_oswt(din_8_rsc_req_obj_oswt),
      .din_8_rsc_req_obj_vd(din_8_rsc_req_obj_vd),
      .din_8_rsc_req_obj_biwt(din_8_rsc_req_obj_biwt),
      .din_8_rsc_req_obj_bdwt(din_8_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj_din_8_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj_din_8_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_8_rsc_req_obj_oswt(din_8_rsc_req_obj_oswt),
      .din_8_rsc_req_obj_wen_comp(din_8_rsc_req_obj_wen_comp),
      .din_8_rsc_req_obj_biwt(din_8_rsc_req_obj_biwt),
      .din_8_rsc_req_obj_bdwt(din_8_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj (
  clk, rst, din_9_rsc_req_vz, core_wen, core_wten, din_9_rsc_req_obj_oswt, din_9_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_9_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_9_rsc_req_obj_oswt;
  output din_9_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_9_rsc_req_obj_vd;
  wire din_9_rsc_req_obj_biwt;
  wire din_9_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_9_rsc_req_obj (
      .vd(din_9_rsc_req_obj_vd),
      .vz(din_9_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj_din_9_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj_din_9_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_9_rsc_req_obj_oswt(din_9_rsc_req_obj_oswt),
      .din_9_rsc_req_obj_vd(din_9_rsc_req_obj_vd),
      .din_9_rsc_req_obj_biwt(din_9_rsc_req_obj_biwt),
      .din_9_rsc_req_obj_bdwt(din_9_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj_din_9_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj_din_9_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_9_rsc_req_obj_oswt(din_9_rsc_req_obj_oswt),
      .din_9_rsc_req_obj_wen_comp(din_9_rsc_req_obj_wen_comp),
      .din_9_rsc_req_obj_biwt(din_9_rsc_req_obj_biwt),
      .din_9_rsc_req_obj_bdwt(din_9_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj (
  clk, rst, din_10_rsc_req_vz, core_wen, core_wten, din_10_rsc_req_obj_oswt, din_10_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_10_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_10_rsc_req_obj_oswt;
  output din_10_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_10_rsc_req_obj_vd;
  wire din_10_rsc_req_obj_biwt;
  wire din_10_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_10_rsc_req_obj (
      .vd(din_10_rsc_req_obj_vd),
      .vz(din_10_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj_din_10_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj_din_10_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_10_rsc_req_obj_oswt(din_10_rsc_req_obj_oswt),
      .din_10_rsc_req_obj_vd(din_10_rsc_req_obj_vd),
      .din_10_rsc_req_obj_biwt(din_10_rsc_req_obj_biwt),
      .din_10_rsc_req_obj_bdwt(din_10_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj_din_10_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj_din_10_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_10_rsc_req_obj_oswt(din_10_rsc_req_obj_oswt),
      .din_10_rsc_req_obj_wen_comp(din_10_rsc_req_obj_wen_comp),
      .din_10_rsc_req_obj_biwt(din_10_rsc_req_obj_biwt),
      .din_10_rsc_req_obj_bdwt(din_10_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj (
  clk, rst, din_11_rsc_req_vz, core_wen, core_wten, din_11_rsc_req_obj_oswt, din_11_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_11_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_11_rsc_req_obj_oswt;
  output din_11_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_11_rsc_req_obj_vd;
  wire din_11_rsc_req_obj_biwt;
  wire din_11_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_11_rsc_req_obj (
      .vd(din_11_rsc_req_obj_vd),
      .vz(din_11_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj_din_11_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj_din_11_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_11_rsc_req_obj_oswt(din_11_rsc_req_obj_oswt),
      .din_11_rsc_req_obj_vd(din_11_rsc_req_obj_vd),
      .din_11_rsc_req_obj_biwt(din_11_rsc_req_obj_biwt),
      .din_11_rsc_req_obj_bdwt(din_11_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj_din_11_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj_din_11_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_11_rsc_req_obj_oswt(din_11_rsc_req_obj_oswt),
      .din_11_rsc_req_obj_wen_comp(din_11_rsc_req_obj_wen_comp),
      .din_11_rsc_req_obj_biwt(din_11_rsc_req_obj_biwt),
      .din_11_rsc_req_obj_bdwt(din_11_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj (
  clk, rst, din_12_rsc_req_vz, core_wen, core_wten, din_12_rsc_req_obj_oswt, din_12_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_12_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_12_rsc_req_obj_oswt;
  output din_12_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_12_rsc_req_obj_vd;
  wire din_12_rsc_req_obj_biwt;
  wire din_12_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_12_rsc_req_obj (
      .vd(din_12_rsc_req_obj_vd),
      .vz(din_12_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj_din_12_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj_din_12_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_12_rsc_req_obj_oswt(din_12_rsc_req_obj_oswt),
      .din_12_rsc_req_obj_vd(din_12_rsc_req_obj_vd),
      .din_12_rsc_req_obj_biwt(din_12_rsc_req_obj_biwt),
      .din_12_rsc_req_obj_bdwt(din_12_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj_din_12_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj_din_12_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_12_rsc_req_obj_oswt(din_12_rsc_req_obj_oswt),
      .din_12_rsc_req_obj_wen_comp(din_12_rsc_req_obj_wen_comp),
      .din_12_rsc_req_obj_biwt(din_12_rsc_req_obj_biwt),
      .din_12_rsc_req_obj_bdwt(din_12_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj (
  clk, rst, din_13_rsc_req_vz, core_wen, core_wten, din_13_rsc_req_obj_oswt, din_13_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_13_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_13_rsc_req_obj_oswt;
  output din_13_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_13_rsc_req_obj_vd;
  wire din_13_rsc_req_obj_biwt;
  wire din_13_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_13_rsc_req_obj (
      .vd(din_13_rsc_req_obj_vd),
      .vz(din_13_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj_din_13_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj_din_13_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_13_rsc_req_obj_oswt(din_13_rsc_req_obj_oswt),
      .din_13_rsc_req_obj_vd(din_13_rsc_req_obj_vd),
      .din_13_rsc_req_obj_biwt(din_13_rsc_req_obj_biwt),
      .din_13_rsc_req_obj_bdwt(din_13_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj_din_13_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj_din_13_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_13_rsc_req_obj_oswt(din_13_rsc_req_obj_oswt),
      .din_13_rsc_req_obj_wen_comp(din_13_rsc_req_obj_wen_comp),
      .din_13_rsc_req_obj_biwt(din_13_rsc_req_obj_biwt),
      .din_13_rsc_req_obj_bdwt(din_13_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj (
  clk, rst, din_14_rsc_req_vz, core_wen, core_wten, din_14_rsc_req_obj_oswt, din_14_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_14_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_14_rsc_req_obj_oswt;
  output din_14_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_14_rsc_req_obj_vd;
  wire din_14_rsc_req_obj_biwt;
  wire din_14_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_14_rsc_req_obj (
      .vd(din_14_rsc_req_obj_vd),
      .vz(din_14_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj_din_14_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj_din_14_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_14_rsc_req_obj_oswt(din_14_rsc_req_obj_oswt),
      .din_14_rsc_req_obj_vd(din_14_rsc_req_obj_vd),
      .din_14_rsc_req_obj_biwt(din_14_rsc_req_obj_biwt),
      .din_14_rsc_req_obj_bdwt(din_14_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj_din_14_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj_din_14_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_14_rsc_req_obj_oswt(din_14_rsc_req_obj_oswt),
      .din_14_rsc_req_obj_wen_comp(din_14_rsc_req_obj_wen_comp),
      .din_14_rsc_req_obj_biwt(din_14_rsc_req_obj_biwt),
      .din_14_rsc_req_obj_bdwt(din_14_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj (
  clk, rst, din_15_rsc_req_vz, core_wen, core_wten, din_15_rsc_req_obj_oswt, din_15_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input din_15_rsc_req_vz;
  input core_wen;
  input core_wten;
  input din_15_rsc_req_obj_oswt;
  output din_15_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_15_rsc_req_obj_vd;
  wire din_15_rsc_req_obj_biwt;
  wire din_15_rsc_req_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v1 #(.valid(32'sd1)) din_15_rsc_req_obj (
      .vd(din_15_rsc_req_obj_vd),
      .vz(din_15_rsc_req_vz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj_din_15_rsc_req_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj_din_15_rsc_req_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_15_rsc_req_obj_oswt(din_15_rsc_req_obj_oswt),
      .din_15_rsc_req_obj_vd(din_15_rsc_req_obj_vd),
      .din_15_rsc_req_obj_biwt(din_15_rsc_req_obj_biwt),
      .din_15_rsc_req_obj_bdwt(din_15_rsc_req_obj_bdwt)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj_din_15_rsc_req_wait_dp
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj_din_15_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_15_rsc_req_obj_oswt(din_15_rsc_req_obj_oswt),
      .din_15_rsc_req_obj_wen_comp(din_15_rsc_req_obj_wen_comp),
      .din_15_rsc_req_obj_biwt(din_15_rsc_req_obj_biwt),
      .din_15_rsc_req_obj_bdwt(din_15_rsc_req_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_rls_obj (
  din_15_rsc_rls_lz, core_wten, din_15_rsc_rls_obj_iswt0
);
  output din_15_rsc_rls_lz;
  input core_wten;
  input din_15_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_15_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_15_rsc_rls_obj (
      .ld(din_15_rsc_rls_obj_ld_core_sct),
      .lz(din_15_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_rls_obj_din_15_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_rls_obj_din_15_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_15_rsc_rls_obj_iswt0(din_15_rsc_rls_obj_iswt0),
      .din_15_rsc_rls_obj_ld_core_sct(din_15_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_rls_obj (
  din_14_rsc_rls_lz, core_wten, din_14_rsc_rls_obj_iswt0
);
  output din_14_rsc_rls_lz;
  input core_wten;
  input din_14_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_14_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_14_rsc_rls_obj (
      .ld(din_14_rsc_rls_obj_ld_core_sct),
      .lz(din_14_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_rls_obj_din_14_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_rls_obj_din_14_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_14_rsc_rls_obj_iswt0(din_14_rsc_rls_obj_iswt0),
      .din_14_rsc_rls_obj_ld_core_sct(din_14_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_rls_obj (
  din_13_rsc_rls_lz, core_wten, din_13_rsc_rls_obj_iswt0
);
  output din_13_rsc_rls_lz;
  input core_wten;
  input din_13_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_13_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_13_rsc_rls_obj (
      .ld(din_13_rsc_rls_obj_ld_core_sct),
      .lz(din_13_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_rls_obj_din_13_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_rls_obj_din_13_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_13_rsc_rls_obj_iswt0(din_13_rsc_rls_obj_iswt0),
      .din_13_rsc_rls_obj_ld_core_sct(din_13_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_rls_obj (
  din_12_rsc_rls_lz, core_wten, din_12_rsc_rls_obj_iswt0
);
  output din_12_rsc_rls_lz;
  input core_wten;
  input din_12_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_12_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_12_rsc_rls_obj (
      .ld(din_12_rsc_rls_obj_ld_core_sct),
      .lz(din_12_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_rls_obj_din_12_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_rls_obj_din_12_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_12_rsc_rls_obj_iswt0(din_12_rsc_rls_obj_iswt0),
      .din_12_rsc_rls_obj_ld_core_sct(din_12_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_rls_obj (
  din_11_rsc_rls_lz, core_wten, din_11_rsc_rls_obj_iswt0
);
  output din_11_rsc_rls_lz;
  input core_wten;
  input din_11_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_11_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_11_rsc_rls_obj (
      .ld(din_11_rsc_rls_obj_ld_core_sct),
      .lz(din_11_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_rls_obj_din_11_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_rls_obj_din_11_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_11_rsc_rls_obj_iswt0(din_11_rsc_rls_obj_iswt0),
      .din_11_rsc_rls_obj_ld_core_sct(din_11_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_rls_obj (
  din_10_rsc_rls_lz, core_wten, din_10_rsc_rls_obj_iswt0
);
  output din_10_rsc_rls_lz;
  input core_wten;
  input din_10_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_10_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_10_rsc_rls_obj (
      .ld(din_10_rsc_rls_obj_ld_core_sct),
      .lz(din_10_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_rls_obj_din_10_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_rls_obj_din_10_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_10_rsc_rls_obj_iswt0(din_10_rsc_rls_obj_iswt0),
      .din_10_rsc_rls_obj_ld_core_sct(din_10_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_rls_obj (
  din_9_rsc_rls_lz, core_wten, din_9_rsc_rls_obj_iswt0
);
  output din_9_rsc_rls_lz;
  input core_wten;
  input din_9_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_9_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_9_rsc_rls_obj (
      .ld(din_9_rsc_rls_obj_ld_core_sct),
      .lz(din_9_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_rls_obj_din_9_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_rls_obj_din_9_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_9_rsc_rls_obj_iswt0(din_9_rsc_rls_obj_iswt0),
      .din_9_rsc_rls_obj_ld_core_sct(din_9_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_rls_obj (
  din_8_rsc_rls_lz, core_wten, din_8_rsc_rls_obj_iswt0
);
  output din_8_rsc_rls_lz;
  input core_wten;
  input din_8_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_8_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_8_rsc_rls_obj (
      .ld(din_8_rsc_rls_obj_ld_core_sct),
      .lz(din_8_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_rls_obj_din_8_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_rls_obj_din_8_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_8_rsc_rls_obj_iswt0(din_8_rsc_rls_obj_iswt0),
      .din_8_rsc_rls_obj_ld_core_sct(din_8_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_rls_obj (
  din_7_rsc_rls_lz, core_wten, din_7_rsc_rls_obj_iswt0
);
  output din_7_rsc_rls_lz;
  input core_wten;
  input din_7_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_7_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_7_rsc_rls_obj (
      .ld(din_7_rsc_rls_obj_ld_core_sct),
      .lz(din_7_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_rls_obj_din_7_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_rls_obj_din_7_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_7_rsc_rls_obj_iswt0(din_7_rsc_rls_obj_iswt0),
      .din_7_rsc_rls_obj_ld_core_sct(din_7_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_rls_obj (
  din_6_rsc_rls_lz, core_wten, din_6_rsc_rls_obj_iswt0
);
  output din_6_rsc_rls_lz;
  input core_wten;
  input din_6_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_6_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_6_rsc_rls_obj (
      .ld(din_6_rsc_rls_obj_ld_core_sct),
      .lz(din_6_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_rls_obj_din_6_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_rls_obj_din_6_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_6_rsc_rls_obj_iswt0(din_6_rsc_rls_obj_iswt0),
      .din_6_rsc_rls_obj_ld_core_sct(din_6_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_rls_obj (
  din_5_rsc_rls_lz, core_wten, din_5_rsc_rls_obj_iswt0
);
  output din_5_rsc_rls_lz;
  input core_wten;
  input din_5_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_5_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_5_rsc_rls_obj (
      .ld(din_5_rsc_rls_obj_ld_core_sct),
      .lz(din_5_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_rls_obj_din_5_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_rls_obj_din_5_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_5_rsc_rls_obj_iswt0(din_5_rsc_rls_obj_iswt0),
      .din_5_rsc_rls_obj_ld_core_sct(din_5_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_rls_obj (
  din_4_rsc_rls_lz, core_wten, din_4_rsc_rls_obj_iswt0
);
  output din_4_rsc_rls_lz;
  input core_wten;
  input din_4_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_4_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_4_rsc_rls_obj (
      .ld(din_4_rsc_rls_obj_ld_core_sct),
      .lz(din_4_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_rls_obj_din_4_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_rls_obj_din_4_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_4_rsc_rls_obj_iswt0(din_4_rsc_rls_obj_iswt0),
      .din_4_rsc_rls_obj_ld_core_sct(din_4_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_rls_obj (
  din_3_rsc_rls_lz, core_wten, din_3_rsc_rls_obj_iswt0
);
  output din_3_rsc_rls_lz;
  input core_wten;
  input din_3_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_3_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_3_rsc_rls_obj (
      .ld(din_3_rsc_rls_obj_ld_core_sct),
      .lz(din_3_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_rls_obj_din_3_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_rls_obj_din_3_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_3_rsc_rls_obj_iswt0(din_3_rsc_rls_obj_iswt0),
      .din_3_rsc_rls_obj_ld_core_sct(din_3_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_rls_obj (
  din_2_rsc_rls_lz, core_wten, din_2_rsc_rls_obj_iswt0
);
  output din_2_rsc_rls_lz;
  input core_wten;
  input din_2_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_2_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_2_rsc_rls_obj (
      .ld(din_2_rsc_rls_obj_ld_core_sct),
      .lz(din_2_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_rls_obj_din_2_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_rls_obj_din_2_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_2_rsc_rls_obj_iswt0(din_2_rsc_rls_obj_iswt0),
      .din_2_rsc_rls_obj_ld_core_sct(din_2_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_rls_obj (
  din_1_rsc_rls_lz, core_wten, din_1_rsc_rls_obj_iswt0
);
  output din_1_rsc_rls_lz;
  input core_wten;
  input din_1_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_1_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_1_rsc_rls_obj (
      .ld(din_1_rsc_rls_obj_ld_core_sct),
      .lz(din_1_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_rls_obj_din_1_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_rls_obj_din_1_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_1_rsc_rls_obj_iswt0(din_1_rsc_rls_obj_iswt0),
      .din_1_rsc_rls_obj_ld_core_sct(din_1_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_rls_obj
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_rls_obj (
  din_0_rsc_rls_lz, core_wten, din_0_rsc_rls_obj_iswt0
);
  output din_0_rsc_rls_lz;
  input core_wten;
  input din_0_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_0_rsc_rls_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v1 #(.valid(32'sd0)) din_0_rsc_rls_obj (
      .ld(din_0_rsc_rls_obj_ld_core_sct),
      .lz(din_0_rsc_rls_lz)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_rls_obj_din_0_rsc_rls_wait_ctrl
      READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_rls_obj_din_0_rsc_rls_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .din_0_rsc_rls_obj_iswt0(din_0_rsc_rls_obj_iswt0),
      .din_0_rsc_rls_obj_ld_core_sct(din_0_rsc_rls_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci (
  clk, rst, dout_rsc_z, dout_rsc_vz, dout_rsc_lz, core_wen, core_wten, dout_rsci_oswt,
      dout_rsci_wen_comp, dout_rsci_d
);
  input clk;
  input rst;
  output [1023:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;
  input core_wen;
  input core_wten;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input [1023:0] dout_rsci_d;


  // Interconnect Declarations
  wire dout_rsci_biwt;
  wire dout_rsci_bdwt;
  wire dout_rsci_ld_core_sct;
  wire dout_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  mgc_out_stdreg_wait_v1 #(.rscid(32'sd161),
  .width(32'sd1024)) dout_rsci (
      .ld(dout_rsci_ld_core_sct),
      .vd(dout_rsci_vd),
      .d(dout_rsci_d),
      .lz(dout_rsc_lz),
      .vz(dout_rsc_vz),
      .z(dout_rsc_z)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_dout_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_dout_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_ld_core_sct(dout_rsci_ld_core_sct),
      .dout_rsci_vd(dout_rsci_vd)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_dout_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_dout_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1 (
  clk, rst, din_15_rsci_douta_d, din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_15_rsci_oswt, din_15_rsci_douta_d_mxwt, din_15_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_15_rsci_douta_d;
  output din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_15_rsci_oswt;
  output [63:0] din_15_rsci_douta_d_mxwt;
  input din_15_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_15_rsci_biwt;
  wire din_15_rsci_bdwt;
  wire din_15_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_din_15_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_din_15_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_15_rsci_oswt(din_15_rsci_oswt),
      .din_15_rsci_biwt(din_15_rsci_biwt),
      .din_15_rsci_bdwt(din_15_rsci_bdwt),
      .din_15_rsci_biwt_pff(din_15_rsci_biwt_iff),
      .din_15_rsci_oswt_pff(din_15_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_din_15_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_din_15_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_15_rsci_douta_d(din_15_rsci_douta_d),
      .din_15_rsci_douta_d_mxwt(din_15_rsci_douta_d_mxwt),
      .din_15_rsci_biwt(din_15_rsci_biwt),
      .din_15_rsci_bdwt(din_15_rsci_bdwt)
    );
  assign din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_15_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1 (
  clk, rst, din_14_rsci_douta_d, din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_14_rsci_oswt, din_14_rsci_douta_d_mxwt, din_14_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_14_rsci_douta_d;
  output din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_14_rsci_oswt;
  output [63:0] din_14_rsci_douta_d_mxwt;
  input din_14_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_14_rsci_biwt;
  wire din_14_rsci_bdwt;
  wire din_14_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_din_14_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_din_14_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_14_rsci_oswt(din_14_rsci_oswt),
      .din_14_rsci_biwt(din_14_rsci_biwt),
      .din_14_rsci_bdwt(din_14_rsci_bdwt),
      .din_14_rsci_biwt_pff(din_14_rsci_biwt_iff),
      .din_14_rsci_oswt_pff(din_14_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_din_14_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_din_14_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_14_rsci_douta_d(din_14_rsci_douta_d),
      .din_14_rsci_douta_d_mxwt(din_14_rsci_douta_d_mxwt),
      .din_14_rsci_biwt(din_14_rsci_biwt),
      .din_14_rsci_bdwt(din_14_rsci_bdwt)
    );
  assign din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_14_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1 (
  clk, rst, din_13_rsci_douta_d, din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_13_rsci_oswt, din_13_rsci_douta_d_mxwt, din_13_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_13_rsci_douta_d;
  output din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_13_rsci_oswt;
  output [63:0] din_13_rsci_douta_d_mxwt;
  input din_13_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_13_rsci_biwt;
  wire din_13_rsci_bdwt;
  wire din_13_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_din_13_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_din_13_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_13_rsci_oswt(din_13_rsci_oswt),
      .din_13_rsci_biwt(din_13_rsci_biwt),
      .din_13_rsci_bdwt(din_13_rsci_bdwt),
      .din_13_rsci_biwt_pff(din_13_rsci_biwt_iff),
      .din_13_rsci_oswt_pff(din_13_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_din_13_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_din_13_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_13_rsci_douta_d(din_13_rsci_douta_d),
      .din_13_rsci_douta_d_mxwt(din_13_rsci_douta_d_mxwt),
      .din_13_rsci_biwt(din_13_rsci_biwt),
      .din_13_rsci_bdwt(din_13_rsci_bdwt)
    );
  assign din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_13_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1 (
  clk, rst, din_12_rsci_douta_d, din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_12_rsci_oswt, din_12_rsci_douta_d_mxwt, din_12_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_12_rsci_douta_d;
  output din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_12_rsci_oswt;
  output [63:0] din_12_rsci_douta_d_mxwt;
  input din_12_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_12_rsci_biwt;
  wire din_12_rsci_bdwt;
  wire din_12_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_din_12_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_din_12_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_12_rsci_oswt(din_12_rsci_oswt),
      .din_12_rsci_biwt(din_12_rsci_biwt),
      .din_12_rsci_bdwt(din_12_rsci_bdwt),
      .din_12_rsci_biwt_pff(din_12_rsci_biwt_iff),
      .din_12_rsci_oswt_pff(din_12_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_din_12_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_din_12_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_12_rsci_douta_d(din_12_rsci_douta_d),
      .din_12_rsci_douta_d_mxwt(din_12_rsci_douta_d_mxwt),
      .din_12_rsci_biwt(din_12_rsci_biwt),
      .din_12_rsci_bdwt(din_12_rsci_bdwt)
    );
  assign din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_12_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1 (
  clk, rst, din_11_rsci_douta_d, din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_11_rsci_oswt, din_11_rsci_douta_d_mxwt, din_11_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_11_rsci_douta_d;
  output din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_11_rsci_oswt;
  output [63:0] din_11_rsci_douta_d_mxwt;
  input din_11_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_11_rsci_biwt;
  wire din_11_rsci_bdwt;
  wire din_11_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_din_11_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_din_11_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_11_rsci_oswt(din_11_rsci_oswt),
      .din_11_rsci_biwt(din_11_rsci_biwt),
      .din_11_rsci_bdwt(din_11_rsci_bdwt),
      .din_11_rsci_biwt_pff(din_11_rsci_biwt_iff),
      .din_11_rsci_oswt_pff(din_11_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_din_11_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_din_11_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_11_rsci_douta_d(din_11_rsci_douta_d),
      .din_11_rsci_douta_d_mxwt(din_11_rsci_douta_d_mxwt),
      .din_11_rsci_biwt(din_11_rsci_biwt),
      .din_11_rsci_bdwt(din_11_rsci_bdwt)
    );
  assign din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_11_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1 (
  clk, rst, din_10_rsci_douta_d, din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, din_10_rsci_oswt, din_10_rsci_douta_d_mxwt, din_10_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_10_rsci_douta_d;
  output din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_10_rsci_oswt;
  output [63:0] din_10_rsci_douta_d_mxwt;
  input din_10_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_10_rsci_biwt;
  wire din_10_rsci_bdwt;
  wire din_10_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_din_10_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_din_10_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_10_rsci_oswt(din_10_rsci_oswt),
      .din_10_rsci_biwt(din_10_rsci_biwt),
      .din_10_rsci_bdwt(din_10_rsci_bdwt),
      .din_10_rsci_biwt_pff(din_10_rsci_biwt_iff),
      .din_10_rsci_oswt_pff(din_10_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_din_10_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_din_10_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_10_rsci_douta_d(din_10_rsci_douta_d),
      .din_10_rsci_douta_d_mxwt(din_10_rsci_douta_d_mxwt),
      .din_10_rsci_biwt(din_10_rsci_biwt),
      .din_10_rsci_bdwt(din_10_rsci_bdwt)
    );
  assign din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_10_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1 (
  clk, rst, din_9_rsci_douta_d, din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_9_rsci_oswt, din_9_rsci_douta_d_mxwt, din_9_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_9_rsci_douta_d;
  output din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_9_rsci_oswt;
  output [63:0] din_9_rsci_douta_d_mxwt;
  input din_9_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_9_rsci_biwt;
  wire din_9_rsci_bdwt;
  wire din_9_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_din_9_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_din_9_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_9_rsci_oswt(din_9_rsci_oswt),
      .din_9_rsci_biwt(din_9_rsci_biwt),
      .din_9_rsci_bdwt(din_9_rsci_bdwt),
      .din_9_rsci_biwt_pff(din_9_rsci_biwt_iff),
      .din_9_rsci_oswt_pff(din_9_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_din_9_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_din_9_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_9_rsci_douta_d(din_9_rsci_douta_d),
      .din_9_rsci_douta_d_mxwt(din_9_rsci_douta_d_mxwt),
      .din_9_rsci_biwt(din_9_rsci_biwt),
      .din_9_rsci_bdwt(din_9_rsci_bdwt)
    );
  assign din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_9_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1 (
  clk, rst, din_8_rsci_douta_d, din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_8_rsci_oswt, din_8_rsci_douta_d_mxwt, din_8_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_8_rsci_douta_d;
  output din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_8_rsci_oswt;
  output [63:0] din_8_rsci_douta_d_mxwt;
  input din_8_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_8_rsci_biwt;
  wire din_8_rsci_bdwt;
  wire din_8_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_din_8_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_din_8_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_8_rsci_oswt(din_8_rsci_oswt),
      .din_8_rsci_biwt(din_8_rsci_biwt),
      .din_8_rsci_bdwt(din_8_rsci_bdwt),
      .din_8_rsci_biwt_pff(din_8_rsci_biwt_iff),
      .din_8_rsci_oswt_pff(din_8_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_din_8_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_din_8_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_8_rsci_douta_d(din_8_rsci_douta_d),
      .din_8_rsci_douta_d_mxwt(din_8_rsci_douta_d_mxwt),
      .din_8_rsci_biwt(din_8_rsci_biwt),
      .din_8_rsci_bdwt(din_8_rsci_bdwt)
    );
  assign din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_8_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1 (
  clk, rst, din_7_rsci_douta_d, din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_7_rsci_oswt, din_7_rsci_douta_d_mxwt, din_7_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_7_rsci_douta_d;
  output din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_7_rsci_oswt;
  output [63:0] din_7_rsci_douta_d_mxwt;
  input din_7_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_7_rsci_biwt;
  wire din_7_rsci_bdwt;
  wire din_7_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_din_7_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_din_7_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_7_rsci_oswt(din_7_rsci_oswt),
      .din_7_rsci_biwt(din_7_rsci_biwt),
      .din_7_rsci_bdwt(din_7_rsci_bdwt),
      .din_7_rsci_biwt_pff(din_7_rsci_biwt_iff),
      .din_7_rsci_oswt_pff(din_7_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_din_7_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_din_7_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_7_rsci_douta_d(din_7_rsci_douta_d),
      .din_7_rsci_douta_d_mxwt(din_7_rsci_douta_d_mxwt),
      .din_7_rsci_biwt(din_7_rsci_biwt),
      .din_7_rsci_bdwt(din_7_rsci_bdwt)
    );
  assign din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_7_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1 (
  clk, rst, din_6_rsci_douta_d, din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_6_rsci_oswt, din_6_rsci_douta_d_mxwt, din_6_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_6_rsci_douta_d;
  output din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_6_rsci_oswt;
  output [63:0] din_6_rsci_douta_d_mxwt;
  input din_6_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_6_rsci_biwt;
  wire din_6_rsci_bdwt;
  wire din_6_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_din_6_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_din_6_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_6_rsci_oswt(din_6_rsci_oswt),
      .din_6_rsci_biwt(din_6_rsci_biwt),
      .din_6_rsci_bdwt(din_6_rsci_bdwt),
      .din_6_rsci_biwt_pff(din_6_rsci_biwt_iff),
      .din_6_rsci_oswt_pff(din_6_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_din_6_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_din_6_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_6_rsci_douta_d(din_6_rsci_douta_d),
      .din_6_rsci_douta_d_mxwt(din_6_rsci_douta_d_mxwt),
      .din_6_rsci_biwt(din_6_rsci_biwt),
      .din_6_rsci_bdwt(din_6_rsci_bdwt)
    );
  assign din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_6_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1 (
  clk, rst, din_5_rsci_douta_d, din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_5_rsci_oswt, din_5_rsci_douta_d_mxwt, din_5_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_5_rsci_douta_d;
  output din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_5_rsci_oswt;
  output [63:0] din_5_rsci_douta_d_mxwt;
  input din_5_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_5_rsci_biwt;
  wire din_5_rsci_bdwt;
  wire din_5_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_din_5_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_din_5_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_5_rsci_oswt(din_5_rsci_oswt),
      .din_5_rsci_biwt(din_5_rsci_biwt),
      .din_5_rsci_bdwt(din_5_rsci_bdwt),
      .din_5_rsci_biwt_pff(din_5_rsci_biwt_iff),
      .din_5_rsci_oswt_pff(din_5_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_din_5_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_din_5_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_5_rsci_douta_d(din_5_rsci_douta_d),
      .din_5_rsci_douta_d_mxwt(din_5_rsci_douta_d_mxwt),
      .din_5_rsci_biwt(din_5_rsci_biwt),
      .din_5_rsci_bdwt(din_5_rsci_bdwt)
    );
  assign din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_5_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1 (
  clk, rst, din_4_rsci_douta_d, din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_4_rsci_oswt, din_4_rsci_douta_d_mxwt, din_4_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_4_rsci_douta_d;
  output din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_4_rsci_oswt;
  output [63:0] din_4_rsci_douta_d_mxwt;
  input din_4_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_4_rsci_biwt;
  wire din_4_rsci_bdwt;
  wire din_4_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_din_4_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_din_4_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_4_rsci_oswt(din_4_rsci_oswt),
      .din_4_rsci_biwt(din_4_rsci_biwt),
      .din_4_rsci_bdwt(din_4_rsci_bdwt),
      .din_4_rsci_biwt_pff(din_4_rsci_biwt_iff),
      .din_4_rsci_oswt_pff(din_4_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_din_4_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_din_4_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_4_rsci_douta_d(din_4_rsci_douta_d),
      .din_4_rsci_douta_d_mxwt(din_4_rsci_douta_d_mxwt),
      .din_4_rsci_biwt(din_4_rsci_biwt),
      .din_4_rsci_bdwt(din_4_rsci_bdwt)
    );
  assign din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_4_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1 (
  clk, rst, din_3_rsci_douta_d, din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_3_rsci_oswt, din_3_rsci_douta_d_mxwt, din_3_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_3_rsci_douta_d;
  output din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_3_rsci_oswt;
  output [63:0] din_3_rsci_douta_d_mxwt;
  input din_3_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_3_rsci_biwt;
  wire din_3_rsci_bdwt;
  wire din_3_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_din_3_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_din_3_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_3_rsci_oswt(din_3_rsci_oswt),
      .din_3_rsci_biwt(din_3_rsci_biwt),
      .din_3_rsci_bdwt(din_3_rsci_bdwt),
      .din_3_rsci_biwt_pff(din_3_rsci_biwt_iff),
      .din_3_rsci_oswt_pff(din_3_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_din_3_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_din_3_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_3_rsci_douta_d(din_3_rsci_douta_d),
      .din_3_rsci_douta_d_mxwt(din_3_rsci_douta_d_mxwt),
      .din_3_rsci_biwt(din_3_rsci_biwt),
      .din_3_rsci_bdwt(din_3_rsci_bdwt)
    );
  assign din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_3_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1 (
  clk, rst, din_2_rsci_douta_d, din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_2_rsci_oswt, din_2_rsci_douta_d_mxwt, din_2_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_2_rsci_douta_d;
  output din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_2_rsci_oswt;
  output [63:0] din_2_rsci_douta_d_mxwt;
  input din_2_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_2_rsci_biwt;
  wire din_2_rsci_bdwt;
  wire din_2_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_din_2_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_din_2_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_2_rsci_oswt(din_2_rsci_oswt),
      .din_2_rsci_biwt(din_2_rsci_biwt),
      .din_2_rsci_bdwt(din_2_rsci_bdwt),
      .din_2_rsci_biwt_pff(din_2_rsci_biwt_iff),
      .din_2_rsci_oswt_pff(din_2_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_din_2_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_din_2_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_2_rsci_douta_d(din_2_rsci_douta_d),
      .din_2_rsci_douta_d_mxwt(din_2_rsci_douta_d_mxwt),
      .din_2_rsci_biwt(din_2_rsci_biwt),
      .din_2_rsci_bdwt(din_2_rsci_bdwt)
    );
  assign din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_2_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1 (
  clk, rst, din_1_rsci_douta_d, din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      core_wten, din_1_rsci_oswt, din_1_rsci_douta_d_mxwt, din_1_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_1_rsci_douta_d;
  output din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input din_1_rsci_oswt;
  output [63:0] din_1_rsci_douta_d_mxwt;
  input din_1_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_1_rsci_biwt;
  wire din_1_rsci_bdwt;
  wire din_1_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_din_1_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_din_1_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_1_rsci_oswt(din_1_rsci_oswt),
      .din_1_rsci_biwt(din_1_rsci_biwt),
      .din_1_rsci_bdwt(din_1_rsci_bdwt),
      .din_1_rsci_biwt_pff(din_1_rsci_biwt_iff),
      .din_1_rsci_oswt_pff(din_1_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_din_1_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_din_1_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_1_rsci_douta_d(din_1_rsci_douta_d),
      .din_1_rsci_douta_d_mxwt(din_1_rsci_douta_d_mxwt),
      .din_1_rsci_biwt(din_1_rsci_biwt),
      .din_1_rsci_bdwt(din_1_rsci_bdwt)
    );
  assign din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_1_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1 (
  clk, rst, din_0_rsci_douta_d, din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, core_wen,
      din_0_rsci_oswt, din_0_rsci_douta_d_mxwt, core_wten, din_0_rsci_oswt_pff
);
  input clk;
  input rst;
  input [63:0] din_0_rsci_douta_d;
  output din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input din_0_rsci_oswt;
  output [63:0] din_0_rsci_douta_d_mxwt;
  input core_wten;
  input din_0_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_0_rsci_biwt;
  wire din_0_rsci_bdwt;
  wire din_0_rsci_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_din_0_rsc_wait_ctrl READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_din_0_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .din_0_rsci_oswt(din_0_rsci_oswt),
      .core_wten(core_wten),
      .din_0_rsci_biwt(din_0_rsci_biwt),
      .din_0_rsci_bdwt(din_0_rsci_bdwt),
      .din_0_rsci_biwt_pff(din_0_rsci_biwt_iff),
      .din_0_rsci_oswt_pff(din_0_rsci_oswt_pff)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_din_0_rsc_wait_dp READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_din_0_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .din_0_rsci_douta_d(din_0_rsci_douta_d),
      .din_0_rsci_douta_d_mxwt(din_0_rsci_douta_d_mxwt),
      .din_0_rsci_biwt(din_0_rsci_biwt),
      .din_0_rsci_bdwt(din_0_rsci_bdwt)
    );
  assign din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_0_rsci_biwt_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, dout_0_rsc_req_vz, dout_0_rsc_rls_lz,
      dout_1_rsc_req_vz, dout_1_rsc_rls_lz, dout_2_rsc_req_vz, dout_2_rsc_rls_lz,
      dout_3_rsc_req_vz, dout_3_rsc_rls_lz, dout_4_rsc_req_vz, dout_4_rsc_rls_lz,
      dout_5_rsc_req_vz, dout_5_rsc_rls_lz, dout_6_rsc_req_vz, dout_6_rsc_rls_lz,
      dout_7_rsc_req_vz, dout_7_rsc_rls_lz, dout_8_rsc_req_vz, dout_8_rsc_rls_lz,
      dout_9_rsc_req_vz, dout_9_rsc_rls_lz, dout_10_rsc_req_vz, dout_10_rsc_rls_lz,
      dout_11_rsc_req_vz, dout_11_rsc_rls_lz, dout_12_rsc_req_vz, dout_12_rsc_rls_lz,
      dout_13_rsc_req_vz, dout_13_rsc_rls_lz, dout_14_rsc_req_vz, dout_14_rsc_rls_lz,
      dout_15_rsc_req_vz, dout_15_rsc_rls_lz, dout_16_rsc_req_vz, dout_16_rsc_rls_lz,
      dout_17_rsc_req_vz, dout_17_rsc_rls_lz, dout_0_rsci_dinb_d, dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_1_rsci_dinb_d, dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_2_rsci_dinb_d,
      dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_3_rsci_dinb_d, dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_4_rsci_dinb_d, dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_5_rsci_dinb_d,
      dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_6_rsci_dinb_d, dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_7_rsci_dinb_d, dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_8_rsci_dinb_d,
      dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_9_rsci_dinb_d, dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_10_rsci_dinb_d, dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_11_rsci_dinb_d,
      dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_12_rsci_dinb_d, dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_13_rsci_dinb_d, dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_14_rsci_dinb_d,
      dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_15_rsci_dinb_d, dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_16_rsci_dinb_d, dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_17_rsci_dinb_d,
      dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_0_data_rsci_addra_d,
      tmp_0_data_rsci_addrb_d, tmp_0_data_rsci_dinb_d, tmp_0_data_rsci_douta_d, tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_1_data_rsci_addra_d,
      tmp_1_data_rsci_addrb_d, tmp_1_data_rsci_dinb_d, tmp_1_data_rsci_douta_d, tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_2_data_rsci_addra_d,
      tmp_2_data_rsci_addrb_d, tmp_2_data_rsci_dinb_d, tmp_2_data_rsci_douta_d, tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_3_data_rsci_addra_d,
      tmp_3_data_rsci_addrb_d, tmp_3_data_rsci_dinb_d, tmp_3_data_rsci_douta_d, tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_4_data_rsci_addra_d,
      tmp_4_data_rsci_addrb_d, tmp_4_data_rsci_dinb_d, tmp_4_data_rsci_douta_d, tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_5_data_rsci_addra_d,
      tmp_5_data_rsci_addrb_d, tmp_5_data_rsci_dinb_d, tmp_5_data_rsci_douta_d, tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_6_data_rsci_addra_d,
      tmp_6_data_rsci_addrb_d, tmp_6_data_rsci_dinb_d, tmp_6_data_rsci_douta_d, tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_7_data_rsci_addra_d,
      tmp_7_data_rsci_addrb_d, tmp_7_data_rsci_dinb_d, tmp_7_data_rsci_douta_d, tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_8_data_rsci_addra_d,
      tmp_8_data_rsci_addrb_d, tmp_8_data_rsci_dinb_d, tmp_8_data_rsci_douta_d, tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_9_data_rsci_addra_d,
      tmp_9_data_rsci_addrb_d, tmp_9_data_rsci_dinb_d, tmp_9_data_rsci_douta_d, tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_10_data_rsci_addra_d,
      tmp_10_data_rsci_addrb_d, tmp_10_data_rsci_dinb_d, tmp_10_data_rsci_douta_d,
      tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      tmp_11_data_rsci_addra_d, tmp_11_data_rsci_addrb_d, tmp_11_data_rsci_dinb_d,
      tmp_11_data_rsci_douta_d, tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_12_data_rsci_addra_d,
      tmp_12_data_rsci_addrb_d, tmp_12_data_rsci_dinb_d, tmp_12_data_rsci_douta_d,
      tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      tmp_13_data_rsci_addra_d, tmp_13_data_rsci_addrb_d, tmp_13_data_rsci_dinb_d,
      tmp_13_data_rsci_douta_d, tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_14_data_rsci_addra_d,
      tmp_14_data_rsci_addrb_d, tmp_14_data_rsci_dinb_d, tmp_14_data_rsci_douta_d,
      tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      tmp_15_data_rsci_addra_d, tmp_15_data_rsci_addrb_d, tmp_15_data_rsci_dinb_d,
      tmp_15_data_rsci_douta_d, tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, tmp_16_data_rsci_addra_d,
      tmp_16_data_rsci_addrb_d, tmp_16_data_rsci_dinb_d, tmp_16_data_rsci_douta_d,
      tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      tmp_17_data_rsci_addra_d, tmp_17_data_rsci_addrb_d, tmp_17_data_rsci_dinb_d,
      tmp_17_data_rsci_douta_d, tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_0_rsci_addra_d_pff,
      dout_1_rsci_addra_d_pff, dout_2_rsci_addra_d_pff, dout_3_rsci_addra_d_pff,
      dout_4_rsci_addra_d_pff, dout_5_rsci_addra_d_pff, dout_6_rsci_addra_d_pff,
      dout_7_rsci_addra_d_pff, dout_8_rsci_addra_d_pff, dout_9_rsci_addra_d_pff,
      dout_10_rsci_addra_d_pff, dout_11_rsci_addra_d_pff, dout_12_rsci_addra_d_pff,
      dout_13_rsci_addra_d_pff, dout_14_rsci_addra_d_pff, dout_15_rsci_addra_d_pff,
      dout_16_rsci_addra_d_pff, dout_17_rsci_addra_d_pff
);
  input clk;
  input rst;
  input [15:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  input dout_0_rsc_req_vz;
  output dout_0_rsc_rls_lz;
  input dout_1_rsc_req_vz;
  output dout_1_rsc_rls_lz;
  input dout_2_rsc_req_vz;
  output dout_2_rsc_rls_lz;
  input dout_3_rsc_req_vz;
  output dout_3_rsc_rls_lz;
  input dout_4_rsc_req_vz;
  output dout_4_rsc_rls_lz;
  input dout_5_rsc_req_vz;
  output dout_5_rsc_rls_lz;
  input dout_6_rsc_req_vz;
  output dout_6_rsc_rls_lz;
  input dout_7_rsc_req_vz;
  output dout_7_rsc_rls_lz;
  input dout_8_rsc_req_vz;
  output dout_8_rsc_rls_lz;
  input dout_9_rsc_req_vz;
  output dout_9_rsc_rls_lz;
  input dout_10_rsc_req_vz;
  output dout_10_rsc_rls_lz;
  input dout_11_rsc_req_vz;
  output dout_11_rsc_rls_lz;
  input dout_12_rsc_req_vz;
  output dout_12_rsc_rls_lz;
  input dout_13_rsc_req_vz;
  output dout_13_rsc_rls_lz;
  input dout_14_rsc_req_vz;
  output dout_14_rsc_rls_lz;
  input dout_15_rsc_req_vz;
  output dout_15_rsc_rls_lz;
  input dout_16_rsc_req_vz;
  output dout_16_rsc_rls_lz;
  input dout_17_rsc_req_vz;
  output dout_17_rsc_rls_lz;
  output [63:0] dout_0_rsci_dinb_d;
  output dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_1_rsci_dinb_d;
  output dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_2_rsci_dinb_d;
  output dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_3_rsci_dinb_d;
  output dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_4_rsci_dinb_d;
  output dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_5_rsci_dinb_d;
  output dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_6_rsci_dinb_d;
  output dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_7_rsci_dinb_d;
  output dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_8_rsci_dinb_d;
  output dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_9_rsci_dinb_d;
  output dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_10_rsci_dinb_d;
  output dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_11_rsci_dinb_d;
  output dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_12_rsci_dinb_d;
  output dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_13_rsci_dinb_d;
  output dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_14_rsci_dinb_d;
  output dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_15_rsci_dinb_d;
  output dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_16_rsci_dinb_d;
  output dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [63:0] dout_17_rsci_dinb_d;
  output dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_0_data_rsci_addra_d;
  output [7:0] tmp_0_data_rsci_addrb_d;
  output [63:0] tmp_0_data_rsci_dinb_d;
  input [63:0] tmp_0_data_rsci_douta_d;
  output tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_1_data_rsci_addra_d;
  output [7:0] tmp_1_data_rsci_addrb_d;
  output [63:0] tmp_1_data_rsci_dinb_d;
  input [63:0] tmp_1_data_rsci_douta_d;
  output tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_2_data_rsci_addra_d;
  output [7:0] tmp_2_data_rsci_addrb_d;
  output [63:0] tmp_2_data_rsci_dinb_d;
  input [63:0] tmp_2_data_rsci_douta_d;
  output tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_3_data_rsci_addra_d;
  output [7:0] tmp_3_data_rsci_addrb_d;
  output [63:0] tmp_3_data_rsci_dinb_d;
  input [63:0] tmp_3_data_rsci_douta_d;
  output tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_4_data_rsci_addra_d;
  output [7:0] tmp_4_data_rsci_addrb_d;
  output [63:0] tmp_4_data_rsci_dinb_d;
  input [63:0] tmp_4_data_rsci_douta_d;
  output tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_5_data_rsci_addra_d;
  output [7:0] tmp_5_data_rsci_addrb_d;
  output [63:0] tmp_5_data_rsci_dinb_d;
  input [63:0] tmp_5_data_rsci_douta_d;
  output tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_6_data_rsci_addra_d;
  output [7:0] tmp_6_data_rsci_addrb_d;
  output [63:0] tmp_6_data_rsci_dinb_d;
  input [63:0] tmp_6_data_rsci_douta_d;
  output tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_7_data_rsci_addra_d;
  output [7:0] tmp_7_data_rsci_addrb_d;
  output [63:0] tmp_7_data_rsci_dinb_d;
  input [63:0] tmp_7_data_rsci_douta_d;
  output tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_8_data_rsci_addra_d;
  output [7:0] tmp_8_data_rsci_addrb_d;
  output [63:0] tmp_8_data_rsci_dinb_d;
  input [63:0] tmp_8_data_rsci_douta_d;
  output tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_9_data_rsci_addra_d;
  output [7:0] tmp_9_data_rsci_addrb_d;
  output [63:0] tmp_9_data_rsci_dinb_d;
  input [63:0] tmp_9_data_rsci_douta_d;
  output tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_10_data_rsci_addra_d;
  output [7:0] tmp_10_data_rsci_addrb_d;
  output [63:0] tmp_10_data_rsci_dinb_d;
  input [63:0] tmp_10_data_rsci_douta_d;
  output tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_11_data_rsci_addra_d;
  output [7:0] tmp_11_data_rsci_addrb_d;
  output [63:0] tmp_11_data_rsci_dinb_d;
  input [63:0] tmp_11_data_rsci_douta_d;
  output tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_12_data_rsci_addra_d;
  output [7:0] tmp_12_data_rsci_addrb_d;
  output [63:0] tmp_12_data_rsci_dinb_d;
  input [63:0] tmp_12_data_rsci_douta_d;
  output tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_13_data_rsci_addra_d;
  output [7:0] tmp_13_data_rsci_addrb_d;
  output [63:0] tmp_13_data_rsci_dinb_d;
  input [63:0] tmp_13_data_rsci_douta_d;
  output tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_14_data_rsci_addra_d;
  output [7:0] tmp_14_data_rsci_addrb_d;
  output [63:0] tmp_14_data_rsci_dinb_d;
  input [63:0] tmp_14_data_rsci_douta_d;
  output tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_15_data_rsci_addra_d;
  output [7:0] tmp_15_data_rsci_addrb_d;
  output [63:0] tmp_15_data_rsci_dinb_d;
  input [63:0] tmp_15_data_rsci_douta_d;
  output tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_16_data_rsci_addra_d;
  output [7:0] tmp_16_data_rsci_addrb_d;
  output [63:0] tmp_16_data_rsci_dinb_d;
  input [63:0] tmp_16_data_rsci_douta_d;
  output tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] tmp_17_data_rsci_addra_d;
  output [7:0] tmp_17_data_rsci_addrb_d;
  output [63:0] tmp_17_data_rsci_dinb_d;
  input [63:0] tmp_17_data_rsci_douta_d;
  output tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [6:0] dout_0_rsci_addra_d_pff;
  output [6:0] dout_1_rsci_addra_d_pff;
  output [6:0] dout_2_rsci_addra_d_pff;
  output [6:0] dout_3_rsci_addra_d_pff;
  output [6:0] dout_4_rsci_addra_d_pff;
  output [6:0] dout_5_rsci_addra_d_pff;
  output [6:0] dout_6_rsci_addra_d_pff;
  output [6:0] dout_7_rsci_addra_d_pff;
  output [6:0] dout_8_rsci_addra_d_pff;
  output [6:0] dout_9_rsci_addra_d_pff;
  output [6:0] dout_10_rsci_addra_d_pff;
  output [6:0] dout_11_rsci_addra_d_pff;
  output [6:0] dout_12_rsci_addra_d_pff;
  output [6:0] dout_13_rsci_addra_d_pff;
  output [6:0] dout_14_rsci_addra_d_pff;
  output [6:0] dout_15_rsci_addra_d_pff;
  output [6:0] dout_16_rsci_addra_d_pff;
  output [6:0] dout_17_rsci_addra_d_pff;


  // Interconnect Declarations
  wire core_wen;
  wire din_rsci_wen_comp;
  wire [15:0] din_rsci_d_mxwt;
  wire core_wten;
  wire [15:0] tmp_0_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_1_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_2_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_3_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_4_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_5_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_6_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_7_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_8_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_9_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_10_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_11_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_12_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_13_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_14_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_15_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_16_data_rsci_douta_d_mxwt;
  wire [15:0] tmp_17_data_rsci_douta_d_mxwt;
  wire dout_17_rsc_req_obj_wen_comp;
  wire dout_16_rsc_req_obj_wen_comp;
  wire dout_15_rsc_req_obj_wen_comp;
  wire dout_14_rsc_req_obj_wen_comp;
  wire dout_13_rsc_req_obj_wen_comp;
  wire dout_12_rsc_req_obj_wen_comp;
  wire dout_11_rsc_req_obj_wen_comp;
  wire dout_10_rsc_req_obj_wen_comp;
  wire dout_9_rsc_req_obj_wen_comp;
  wire dout_8_rsc_req_obj_wen_comp;
  wire dout_7_rsc_req_obj_wen_comp;
  wire dout_6_rsc_req_obj_wen_comp;
  wire dout_5_rsc_req_obj_wen_comp;
  wire dout_4_rsc_req_obj_wen_comp;
  wire dout_3_rsc_req_obj_wen_comp;
  wire dout_2_rsc_req_obj_wen_comp;
  wire dout_1_rsc_req_obj_wen_comp;
  wire dout_0_rsc_req_obj_wen_comp;
  wire [4:0] mux1h_77_tmp;
  wire [4:0] mux1h_78_tmp;
  wire or_2_tmp_1;
  wire nor_19_tmp;
  wire [6:0] mux1h_19_tmp;
  wire [6:0] mux1h_18_tmp;
  wire [6:0] mux1h_17_tmp;
  wire [6:0] mux1h_16_tmp;
  wire [6:0] mux1h_15_tmp;
  wire [6:0] mux1h_14_tmp;
  wire [6:0] mux1h_13_tmp;
  wire [6:0] mux1h_12_tmp;
  wire [6:0] mux1h_11_tmp;
  wire [6:0] mux1h_10_tmp;
  wire [6:0] mux1h_9_tmp;
  wire [6:0] mux1h_8_tmp;
  wire [6:0] mux1h_7_tmp;
  wire [6:0] mux1h_6_tmp;
  wire [6:0] mux1h_5_tmp;
  wire [6:0] mux1h_4_tmp;
  wire [6:0] mux1h_3_tmp;
  wire and_dcpl_19;
  wire and_dcpl_20;
  wire or_dcpl_8;
  wire or_dcpl_10;
  wire or_dcpl_11;
  wire or_dcpl_12;
  wire or_dcpl_15;
  wire or_dcpl_16;
  wire or_dcpl_17;
  wire or_dcpl_24;
  wire or_dcpl_28;
  wire or_dcpl_36;
  wire or_dcpl_37;
  wire or_dcpl_38;
  wire or_dcpl_41;
  wire or_dcpl_42;
  wire or_dcpl_43;
  wire or_dcpl_53;
  wire or_dcpl_61;
  wire or_dcpl_80;
  wire or_dcpl_81;
  wire or_dcpl_84;
  wire or_dcpl_101;
  wire or_dcpl_102;
  wire or_dcpl_121;
  wire or_dcpl_124;
  wire or_dcpl_141;
  wire or_dcpl_160;
  wire or_dcpl_161;
  wire or_dcpl_164;
  wire or_dcpl_181;
  wire or_dcpl_194;
  wire or_dcpl_195;
  wire or_dcpl_196;
  wire or_dcpl_197;
  wire or_dcpl_198;
  wire or_dcpl_200;
  wire or_dcpl_201;
  wire or_dcpl_202;
  wire or_dcpl_204;
  wire or_dcpl_205;
  wire or_dcpl_207;
  wire or_dcpl_208;
  wire or_dcpl_210;
  wire or_dcpl_211;
  wire or_dcpl_213;
  wire or_dcpl_214;
  wire or_dcpl_215;
  wire or_dcpl_217;
  wire or_dcpl_218;
  wire or_dcpl_220;
  wire or_dcpl_221;
  wire or_dcpl_223;
  wire or_dcpl_224;
  wire or_dcpl_226;
  wire or_dcpl_228;
  wire or_dcpl_230;
  wire or_dcpl_232;
  wire or_dcpl_233;
  wire or_dcpl_235;
  wire or_dcpl_237;
  wire or_dcpl_239;
  wire or_dcpl_241;
  wire or_dcpl_243;
  wire or_dcpl_246;
  wire or_dcpl_248;
  wire or_dcpl_249;
  wire or_dcpl_250;
  wire or_dcpl_251;
  wire or_dcpl_253;
  wire or_dcpl_256;
  wire or_dcpl_257;
  wire or_dcpl_260;
  wire or_tmp_75;
  wire or_dcpl_262;
  wire or_dcpl_263;
  wire or_dcpl_264;
  wire nor_tmp_21;
  wire or_dcpl_267;
  wire or_dcpl_268;
  wire or_dcpl_271;
  wire or_dcpl_272;
  wire or_dcpl_275;
  wire or_dcpl_277;
  wire or_dcpl_278;
  wire or_dcpl_279;
  wire or_tmp_82;
  wire or_dcpl_281;
  wire nor_tmp_23;
  wire or_dcpl_284;
  wire or_dcpl_286;
  wire or_dcpl_289;
  wire or_dcpl_293;
  wire nor_tmp_25;
  wire or_tmp_90;
  wire mux_tmp_42;
  wire nor_tmp_26;
  wire or_dcpl_302;
  wire or_tmp_101;
  wire nor_tmp_28;
  wire or_dcpl_307;
  wire or_dcpl_312;
  wire and_dcpl_28;
  reg [6:0] WRITE_x_idx_6_0_lpi_2;
  reg lfst_exit_WRITE_lpi_1;
  reg [4:0] WRITE_for_y_idx_4_0_lpi_3;
  reg [6:0] io_write_dout_0_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_1_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_2_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_3_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_4_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_5_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_6_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_7_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_8_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_9_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_10_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_11_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_12_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_13_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_14_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_15_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_16_copy_ndx_6_0_lpi_1;
  reg [6:0] io_write_dout_17_copy_ndx_6_0_lpi_1;
  reg exit_WRITE_sva_2;
  reg [6:0] io_write_dout_17_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_17_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_17_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_16_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_16_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_16_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_15_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_15_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_15_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_14_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_14_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_14_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_13_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_13_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_13_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_12_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_12_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_12_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_11_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_11_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_11_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_10_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_10_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_10_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_9_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_9_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_9_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_8_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_8_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_8_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_7_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_7_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_7_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_6_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_6_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_6_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_5_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_5_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_5_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_4_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_4_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_4_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_3_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_3_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_3_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_2_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_2_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_2_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_1_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_1_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_1_copy_ndx_6_0_lpi_1_dfm_4;
  reg [6:0] io_write_dout_0_copy_ndx_6_0_sva_4;
  wire [7:0] nl_io_write_dout_0_copy_ndx_6_0_sva_4;
  reg [6:0] io_write_dout_0_copy_ndx_6_0_lpi_1_dfm_4;
  reg exit_WRITE_lpi_1_dfm_4;
  reg WRITE_for_slc_WRITE_for_acc_4_svs_2;
  reg [4:0] WRITE_for_y_idx_4_0_sva_6;
  reg [6:0] WRITE_x_idx_6_0_lpi_1_dfm_5;
  reg [4:0] lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24;
  reg equal_tmp_18;
  reg equal_tmp_72;
  reg equal_tmp_20;
  reg equal_tmp_73;
  reg equal_tmp_22;
  reg equal_tmp_74;
  reg equal_tmp_24;
  reg equal_tmp_75;
  reg equal_tmp_26;
  reg equal_tmp_76;
  reg equal_tmp_28;
  reg equal_tmp_77;
  reg equal_tmp_30;
  reg equal_tmp_78;
  reg equal_tmp_32;
  reg equal_tmp_79;
  reg equal_tmp_34;
  reg equal_tmp_80;
  reg equal_tmp_36;
  reg equal_tmp_81;
  reg equal_tmp_38;
  reg equal_tmp_82;
  reg equal_tmp_40;
  reg equal_tmp_83;
  reg equal_tmp_42;
  reg equal_tmp_84;
  reg equal_tmp_44;
  reg equal_tmp_85;
  reg equal_tmp_46;
  reg equal_tmp_86;
  reg equal_tmp_48;
  reg equal_tmp_87;
  reg equal_tmp_50;
  reg equal_tmp_88;
  reg equal_tmp_52;
  reg equal_tmp_89;
  reg nor_tmp_1;
  reg nor_tmp_30;
  reg nor_dfs_3;
  reg [4:0] WRITE_for_y_idx_4_0_lpi_1_dfm_st_2;
  reg WRITE_for_y_idx_slc_WRITE_for_y_idx_4_0_0_itm_3;
  reg [4:0] lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3;
  reg main_stage_0_2;
  reg main_stage_0_3;
  wire lfst_exit_WRITE_lpi_1_mx0;
  wire for_unequal_tmp;
  wire unequal_tmp;
  wire unequal_tmp_1;
  wire unequal_tmp_2;
  wire unequal_tmp_3;
  wire unequal_tmp_4;
  wire unequal_tmp_5;
  wire unequal_tmp_6;
  wire unequal_tmp_7;
  wire unequal_tmp_8;
  wire unequal_tmp_9;
  wire unequal_tmp_10;
  wire unequal_tmp_11;
  wire unequal_tmp_12;
  wire unequal_tmp_13;
  wire unequal_tmp_14;
  wire unequal_tmp_15;
  wire unequal_tmp_16;
  wire equal_tmp;
  wire equal_tmp_1;
  wire equal_tmp_2;
  wire equal_tmp_3;
  wire equal_tmp_4;
  wire equal_tmp_5;
  wire equal_tmp_6;
  wire equal_tmp_7;
  wire equal_tmp_8;
  wire equal_tmp_9;
  wire equal_tmp_10;
  wire equal_tmp_11;
  wire equal_tmp_12;
  wire equal_tmp_13;
  wire equal_tmp_14;
  wire equal_tmp_15;
  wire equal_tmp_16;
  wire equal_tmp_17;
  wire nor_tmp;
  wire [6:0] io_write_dout_0_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_1_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_2_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_3_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_4_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_5_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_6_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_7_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_8_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_9_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_10_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_11_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_12_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_13_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_14_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_15_copy_ndx_6_0_lpi_1_mx0;
  wire [6:0] io_write_dout_16_copy_ndx_6_0_lpi_1_mx0;
  wire [4:0] lfst_exit_io_write_dout_17_copy_lpi_1_dfm;
  wire [6:0] WRITE_x_idx_6_0_sva_1;
  wire [7:0] nl_WRITE_x_idx_6_0_sva_1;
  wire or_3_tmp;
  wire or_4_tmp;
  wire or_5_tmp;
  wire or_6_tmp;
  wire or_7_tmp;
  wire or_8_tmp;
  wire or_9_tmp;
  wire or_10_tmp;
  wire or_11_tmp;
  wire or_12_tmp;
  wire or_13_tmp;
  wire or_14_tmp;
  wire or_15_tmp;
  wire or_16_tmp;
  wire or_17_tmp;
  wire or_18_tmp;
  wire or_19_tmp;
  wire or_20_tmp;
  wire [6:0] mux_53_tmp;
  wire and_76_rgt;
  wire or_1_tmp;
  reg reg_dout_0_rsc_rls_obj_iswt0_cse;
  reg reg_dout_1_rsc_rls_obj_iswt0_cse;
  reg reg_dout_2_rsc_rls_obj_iswt0_cse;
  reg reg_dout_3_rsc_rls_obj_iswt0_cse;
  reg reg_dout_4_rsc_rls_obj_iswt0_cse;
  reg reg_dout_5_rsc_rls_obj_iswt0_cse;
  reg reg_dout_6_rsc_rls_obj_iswt0_cse;
  reg reg_dout_7_rsc_rls_obj_iswt0_cse;
  reg reg_dout_8_rsc_rls_obj_iswt0_cse;
  reg reg_dout_9_rsc_rls_obj_iswt0_cse;
  reg reg_dout_10_rsc_rls_obj_iswt0_cse;
  reg reg_dout_11_rsc_rls_obj_iswt0_cse;
  reg reg_dout_12_rsc_rls_obj_iswt0_cse;
  reg reg_dout_13_rsc_rls_obj_iswt0_cse;
  reg reg_dout_14_rsc_rls_obj_iswt0_cse;
  reg reg_dout_15_rsc_rls_obj_iswt0_cse;
  reg reg_dout_16_rsc_rls_obj_iswt0_cse;
  reg reg_dout_17_rsc_rls_obj_iswt0_cse;
  reg reg_dout_17_rsc_req_obj_oswt_cse;
  reg reg_dout_16_rsc_req_obj_oswt_cse;
  reg reg_dout_15_rsc_req_obj_oswt_cse;
  reg reg_dout_14_rsc_req_obj_oswt_cse;
  reg reg_dout_13_rsc_req_obj_oswt_cse;
  reg reg_dout_12_rsc_req_obj_oswt_cse;
  reg reg_dout_11_rsc_req_obj_oswt_cse;
  reg reg_dout_10_rsc_req_obj_oswt_cse;
  reg reg_dout_9_rsc_req_obj_oswt_cse;
  reg reg_dout_8_rsc_req_obj_oswt_cse;
  reg reg_dout_7_rsc_req_obj_oswt_cse;
  reg reg_dout_6_rsc_req_obj_oswt_cse;
  reg reg_dout_5_rsc_req_obj_oswt_cse;
  reg reg_dout_4_rsc_req_obj_oswt_cse;
  reg reg_dout_3_rsc_req_obj_oswt_cse;
  reg reg_dout_2_rsc_req_obj_oswt_cse;
  reg reg_dout_1_rsc_req_obj_oswt_cse;
  reg reg_tmp_0_data_rsci_oswt_cse;
  reg reg_tmp_1_data_rsci_oswt_cse;
  reg reg_tmp_2_data_rsci_oswt_cse;
  reg reg_tmp_3_data_rsci_oswt_cse;
  reg reg_tmp_4_data_rsci_oswt_cse;
  reg reg_tmp_5_data_rsci_oswt_cse;
  reg reg_tmp_6_data_rsci_oswt_cse;
  reg reg_tmp_7_data_rsci_oswt_cse;
  reg reg_tmp_8_data_rsci_oswt_cse;
  reg reg_tmp_9_data_rsci_oswt_cse;
  reg reg_tmp_10_data_rsci_oswt_cse;
  reg reg_tmp_11_data_rsci_oswt_cse;
  reg reg_tmp_12_data_rsci_oswt_cse;
  reg reg_tmp_13_data_rsci_oswt_cse;
  reg reg_tmp_14_data_rsci_oswt_cse;
  reg reg_tmp_15_data_rsci_oswt_cse;
  reg reg_tmp_16_data_rsci_oswt_cse;
  reg reg_tmp_17_data_rsci_oswt_cse;
  reg reg_dout_0_rsc_req_obj_oswt_cse;
  reg reg_din_rsci_oswt_cse;
  wire [63:0] dout_0_rsci_dinb_d_reg;
  wire dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_1_rsci_dinb_d_reg;
  wire dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_2_rsci_dinb_d_reg;
  wire dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_3_rsci_dinb_d_reg;
  wire dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_4_rsci_dinb_d_reg;
  wire dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_5_rsci_dinb_d_reg;
  wire dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_6_rsci_dinb_d_reg;
  wire dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_7_rsci_dinb_d_reg;
  wire dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_8_rsci_dinb_d_reg;
  wire dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_9_rsci_dinb_d_reg;
  wire dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_10_rsci_dinb_d_reg;
  wire dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_11_rsci_dinb_d_reg;
  wire dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_12_rsci_dinb_d_reg;
  wire dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_13_rsci_dinb_d_reg;
  wire dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_14_rsci_dinb_d_reg;
  wire dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_15_rsci_dinb_d_reg;
  wire dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_16_rsci_dinb_d_reg;
  wire dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [63:0] dout_17_rsci_dinb_d_reg;
  wire dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_0_data_rsci_addra_d_reg;
  wire WRITE_for_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_rmff;
  wire [7:0] tmp_0_data_rsci_addrb_d_reg;
  wire tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_1_data_rsci_addra_d_reg;
  wire WRITE_for_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_1_rmff;
  wire [7:0] tmp_1_data_rsci_addrb_d_reg;
  wire tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_2_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_2_rmff;
  wire [7:0] tmp_2_data_rsci_addrb_d_reg;
  wire tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_3_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_3_rmff;
  wire [7:0] tmp_3_data_rsci_addrb_d_reg;
  wire tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_4_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_4_rmff;
  wire [7:0] tmp_4_data_rsci_addrb_d_reg;
  wire tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_5_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_5_rmff;
  wire [7:0] tmp_5_data_rsci_addrb_d_reg;
  wire tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_6_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_6_rmff;
  wire [7:0] tmp_6_data_rsci_addrb_d_reg;
  wire tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_7_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_7_rmff;
  wire [7:0] tmp_7_data_rsci_addrb_d_reg;
  wire tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_8_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_8_rmff;
  wire [7:0] tmp_8_data_rsci_addrb_d_reg;
  wire tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_9_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_9_rmff;
  wire [7:0] tmp_9_data_rsci_addrb_d_reg;
  wire tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_10_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_10_rmff;
  wire [7:0] tmp_10_data_rsci_addrb_d_reg;
  wire tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_11_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_11_rmff;
  wire [7:0] tmp_11_data_rsci_addrb_d_reg;
  wire tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_12_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_12_rmff;
  wire [7:0] tmp_12_data_rsci_addrb_d_reg;
  wire tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_13_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_13_rmff;
  wire [7:0] tmp_13_data_rsci_addrb_d_reg;
  wire tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_14_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_14_rmff;
  wire [7:0] tmp_14_data_rsci_addrb_d_reg;
  wire tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_15_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_15_rmff;
  wire [7:0] tmp_15_data_rsci_addrb_d_reg;
  wire tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_16_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_16_rmff;
  wire [7:0] tmp_16_data_rsci_addrb_d_reg;
  wire tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [7:0] tmp_17_data_rsci_addra_d_reg;
  wire WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
  wire [6:0] WRITE_x_idx_mux_17_rmff;
  wire [7:0] tmp_17_data_rsci_addrb_d_reg;
  wire tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire or_732_tmp;
  wire nor_tmp_31;
  wire [4:0] WRITE_for_y_idx_4_0_sva_1;
  wire [5:0] nl_WRITE_for_y_idx_4_0_sva_1;
  wire [4:0] WRITE_for_y_idx_4_0_lpi_1_dfm;
  wire [6:0] WRITE_x_idx_6_0_lpi_1_dfm;
  wire and_206_cse;
  wire and_208_cse;
  wire and_210_cse;
  wire and_212_cse;
  wire and_214_cse;
  wire and_216_cse;
  wire and_218_cse;
  wire and_220_cse;
  wire and_222_cse;
  wire and_224_cse;
  wire and_226_cse;
  wire and_228_cse;
  wire and_230_cse;
  wire and_232_cse;
  wire and_234_cse;
  wire and_236_cse;
  wire and_238_cse;
  wire mux_130_cse;
  wire WRITE_for_acc_itm_4_1;
  wire WRITE_acc_itm_6;

  wire[0:0] mux_132_nl;
  wire[0:0] and_141_nl;
  wire[0:0] or_245_nl;
  wire[0:0] nor_76_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] and_142_nl;
  wire[0:0] or_253_nl;
  wire[0:0] nor_77_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] and_143_nl;
  wire[0:0] or_260_nl;
  wire[0:0] nor_78_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] and_144_nl;
  wire[0:0] or_270_nl;
  wire[0:0] nor_79_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] and_145_nl;
  wire[0:0] or_278_nl;
  wire[0:0] nor_80_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] and_146_nl;
  wire[0:0] or_285_nl;
  wire[0:0] nor_81_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] and_147_nl;
  wire[0:0] or_292_nl;
  wire[0:0] nor_82_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] and_148_nl;
  wire[0:0] or_299_nl;
  wire[0:0] nor_83_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] and_149_nl;
  wire[0:0] or_305_nl;
  wire[0:0] nor_84_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] and_150_nl;
  wire[0:0] or_311_nl;
  wire[0:0] nor_85_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] and_151_nl;
  wire[0:0] or_317_nl;
  wire[0:0] nor_86_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] and_152_nl;
  wire[0:0] or_324_nl;
  wire[0:0] nor_87_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] and_153_nl;
  wire[0:0] or_330_nl;
  wire[0:0] nor_88_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] and_154_nl;
  wire[0:0] or_336_nl;
  wire[0:0] nor_89_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] and_155_nl;
  wire[0:0] or_342_nl;
  wire[0:0] nor_90_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] and_156_nl;
  wire[0:0] or_348_nl;
  wire[0:0] nor_91_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] and_157_nl;
  wire[0:0] or_354_nl;
  wire[0:0] nor_92_nl;
  wire[0:0] WRITE_not_8_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] or_358_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] or_359_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] and_168_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] nor_116_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] or_375_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] nor_114_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] or_388_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] nor_113_nl;
  wire[0:0] and_166_nl;
  wire[0:0] mux_164_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] or_400_nl;
  wire[0:0] nor_111_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] or_408_nl;
  wire[0:0] nor_110_nl;
  wire[0:0] mux_168_nl;
  wire[0:0] or_415_nl;
  wire[0:0] mux_167_nl;
  wire[0:0] or_416_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] and_164_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] nor_108_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] or_426_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] nor_107_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] or_433_nl;
  wire[0:0] or_435_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] mux_180_nl;
  wire[0:0] nor_106_nl;
  wire[0:0] and_161_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] or_442_nl;
  wire[0:0] nor_104_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] mux_184_nl;
  wire[0:0] or_449_nl;
  wire[0:0] nor_103_nl;
  wire[0:0] mux_186_nl;
  wire[0:0] or_454_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] nor_102_nl;
  wire[0:0] or_568_nl;
  wire[0:0] and_190_nl;
  wire[0:0] and_191_nl;
  wire[0:0] and_169_nl;
  wire[4:0] WRITE_for_acc_nl;
  wire[5:0] nl_WRITE_for_acc_nl;
  wire[0:0] for_for_and_1_nl;
  wire[0:0] nor_257_nl;
  wire[0:0] or_472_nl;
  wire[1:0] for_mux_3_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] and_202_nl;
  wire[0:0] and_79_nl;
  wire[0:0] and_81_nl;
  wire[0:0] and_83_nl;
  wire[0:0] and_85_nl;
  wire[0:0] and_87_nl;
  wire[0:0] and_89_nl;
  wire[0:0] and_91_nl;
  wire[0:0] and_93_nl;
  wire[0:0] and_95_nl;
  wire[0:0] and_97_nl;
  wire[0:0] and_99_nl;
  wire[0:0] and_101_nl;
  wire[0:0] and_103_nl;
  wire[0:0] and_105_nl;
  wire[0:0] and_107_nl;
  wire[0:0] and_109_nl;
  wire[0:0] and_111_nl;
  wire[0:0] and_203_nl;
  wire[6:0] WRITE_acc_nl;
  wire[7:0] nl_WRITE_acc_nl;
  wire[0:0] nor_117_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_inst_dout_0_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_inst_dout_0_rsci_dinb_d_core
      = {48'b0, tmp_0_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_inst_dout_0_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_inst_dout_0_rsci_iswt0_pff
      = ~(or_dcpl_17 | or_dcpl_16);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_inst_dout_1_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_inst_dout_1_rsci_dinb_d_core
      = {48'b0, tmp_1_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_inst_dout_1_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_inst_dout_1_rsci_iswt0_pff
      = ~(or_dcpl_17 | or_dcpl_28);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_inst_dout_2_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_inst_dout_2_rsci_dinb_d_core
      = {48'b0, tmp_2_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_inst_dout_2_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_inst_dout_2_rsci_iswt0_pff
      = ~(or_dcpl_43 | or_dcpl_42);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_inst_dout_3_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_inst_dout_3_rsci_dinb_d_core
      = {48'b0, tmp_3_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_inst_dout_3_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_inst_dout_3_rsci_iswt0_pff
      = ~(or_dcpl_43 | or_dcpl_53);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_inst_dout_4_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_inst_dout_4_rsci_dinb_d_core
      = {48'b0, tmp_4_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_inst_dout_4_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_inst_dout_4_rsci_iswt0_pff
      = ~(or_dcpl_43 | or_dcpl_16);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_inst_dout_5_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_inst_dout_5_rsci_dinb_d_core
      = {48'b0, tmp_5_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_inst_dout_5_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_inst_dout_5_rsci_iswt0_pff
      = ~(or_dcpl_43 | or_dcpl_28);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_inst_dout_6_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_inst_dout_6_rsci_dinb_d_core
      = {48'b0, tmp_6_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_inst_dout_6_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_inst_dout_6_rsci_iswt0_pff
      = ~(or_dcpl_84 | or_dcpl_42);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_inst_dout_7_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_inst_dout_7_rsci_dinb_d_core
      = {48'b0, tmp_7_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_inst_dout_7_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_inst_dout_7_rsci_iswt0_pff
      = ~(or_dcpl_84 | or_dcpl_53);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_inst_dout_8_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_inst_dout_8_rsci_dinb_d_core
      = {48'b0, tmp_8_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_inst_dout_8_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_inst_dout_8_rsci_iswt0_pff
      = ~(or_dcpl_84 | or_dcpl_16);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_inst_dout_9_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_inst_dout_9_rsci_dinb_d_core
      = {48'b0, tmp_9_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_inst_dout_9_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_inst_dout_9_rsci_iswt0_pff
      = ~(or_dcpl_84 | or_dcpl_28);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_inst_dout_10_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_inst_dout_10_rsci_dinb_d_core
      = {48'b0, tmp_10_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_inst_dout_10_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_inst_dout_10_rsci_iswt0_pff
      = ~(or_dcpl_124 | or_dcpl_42);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_inst_dout_11_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_inst_dout_11_rsci_dinb_d_core
      = {48'b0, tmp_11_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_inst_dout_11_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_inst_dout_11_rsci_iswt0_pff
      = ~(or_dcpl_124 | or_dcpl_53);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_inst_dout_12_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_inst_dout_12_rsci_dinb_d_core
      = {48'b0, tmp_12_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_inst_dout_12_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_inst_dout_12_rsci_iswt0_pff
      = ~(or_dcpl_124 | or_dcpl_16);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_inst_dout_13_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_inst_dout_13_rsci_dinb_d_core
      = {48'b0, tmp_13_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_inst_dout_13_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_inst_dout_13_rsci_iswt0_pff
      = ~(or_dcpl_124 | or_dcpl_28);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_inst_dout_14_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_inst_dout_14_rsci_dinb_d_core
      = {48'b0, tmp_14_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_inst_dout_14_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_inst_dout_14_rsci_iswt0_pff
      = ~(or_dcpl_164 | or_dcpl_42);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_inst_dout_15_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_inst_dout_15_rsci_dinb_d_core
      = {48'b0, tmp_15_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_inst_dout_15_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_inst_dout_15_rsci_iswt0_pff
      = ~(or_dcpl_164 | or_dcpl_53);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_inst_dout_16_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_inst_dout_16_rsci_dinb_d_core
      = {48'b0, tmp_16_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_inst_dout_16_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_inst_dout_16_rsci_iswt0_pff
      = ~(or_dcpl_164 | or_dcpl_16);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [63:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_inst_dout_17_rsci_dinb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_inst_dout_17_rsci_dinb_d_core
      = {48'b0, tmp_17_data_rsci_douta_d_mxwt};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_inst_dout_17_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_inst_dout_17_rsci_iswt0_pff
      = ~(or_dcpl_164 | or_dcpl_28);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_243;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_253 | or_dcpl_251);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_1_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_1_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_241;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_253 | or_dcpl_257);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_2_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_2_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_239;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_253 | or_dcpl_264);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_3_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_3_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_237;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_253 | or_dcpl_268);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_4_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_4_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_235;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_253 | or_dcpl_272);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_5_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_5_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_233;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_253 | or_dcpl_275);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_6_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_6_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_230;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_253 | or_dcpl_281);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_7_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_7_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_228;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_253 | or_dcpl_284);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_8_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_8_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_226;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_289 | or_dcpl_251);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_9_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_9_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_224;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_289 | or_dcpl_257);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_10_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_10_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_221;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_289 | or_dcpl_264);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_11_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_11_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_218;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_289 | or_dcpl_268);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_12_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_12_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_215;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_289 | or_dcpl_272);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_13_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_13_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_211;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_289 | or_dcpl_275);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_14_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_14_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_205;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_289 | or_dcpl_281);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_15_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_15_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_202;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_289 | or_dcpl_284);
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_16_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_16_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~ or_dcpl_198;
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_312 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]) | WRITE_for_y_idx_slc_WRITE_for_y_idx_4_0_0_itm_3
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]));
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_addra_d_core
      = {1'b0, WRITE_x_idx_mux_17_rmff};
  wire [7:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_addrb_d_core
      = {1'b0, WRITE_x_idx_mux_17_rmff};
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct
      = ~(or_dcpl_197 | or_dcpl_223);
  wire [0:0] nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct;
  assign nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct
      = ~(or_dcpl_312 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]) | (~ WRITE_for_y_idx_slc_WRITE_for_y_idx_4_0_0_itm_3)
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]));
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_din_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(din_rsc_z),
      .din_rsc_vz(din_rsc_vz),
      .din_rsc_lz(din_rsc_lz),
      .core_wen(core_wen),
      .din_rsci_oswt(reg_din_rsci_oswt_cse),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_d_mxwt(din_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_inst
      (
      .dout_0_rsci_dinb_d(dout_0_rsci_dinb_d_reg),
      .dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_0_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_inst_dout_0_rsci_dinb_d_core[63:0]),
      .dout_0_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_inst_dout_0_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_inst
      (
      .dout_1_rsci_dinb_d(dout_1_rsci_dinb_d_reg),
      .dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_1_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_inst_dout_1_rsci_dinb_d_core[63:0]),
      .dout_1_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_inst_dout_1_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_inst
      (
      .dout_2_rsci_dinb_d(dout_2_rsci_dinb_d_reg),
      .dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_2_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_inst_dout_2_rsci_dinb_d_core[63:0]),
      .dout_2_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_inst_dout_2_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_inst
      (
      .dout_3_rsci_dinb_d(dout_3_rsci_dinb_d_reg),
      .dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_3_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_inst_dout_3_rsci_dinb_d_core[63:0]),
      .dout_3_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_inst_dout_3_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_inst
      (
      .dout_4_rsci_dinb_d(dout_4_rsci_dinb_d_reg),
      .dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_4_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_inst_dout_4_rsci_dinb_d_core[63:0]),
      .dout_4_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_inst_dout_4_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_inst
      (
      .dout_5_rsci_dinb_d(dout_5_rsci_dinb_d_reg),
      .dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_5_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_inst_dout_5_rsci_dinb_d_core[63:0]),
      .dout_5_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_inst_dout_5_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_inst
      (
      .dout_6_rsci_dinb_d(dout_6_rsci_dinb_d_reg),
      .dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_6_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_inst_dout_6_rsci_dinb_d_core[63:0]),
      .dout_6_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_inst_dout_6_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_inst
      (
      .dout_7_rsci_dinb_d(dout_7_rsci_dinb_d_reg),
      .dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_7_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_inst_dout_7_rsci_dinb_d_core[63:0]),
      .dout_7_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_inst_dout_7_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_inst
      (
      .dout_8_rsci_dinb_d(dout_8_rsci_dinb_d_reg),
      .dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_8_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_inst_dout_8_rsci_dinb_d_core[63:0]),
      .dout_8_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_inst_dout_8_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_inst
      (
      .dout_9_rsci_dinb_d(dout_9_rsci_dinb_d_reg),
      .dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_9_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_inst_dout_9_rsci_dinb_d_core[63:0]),
      .dout_9_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_inst_dout_9_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_inst
      (
      .dout_10_rsci_dinb_d(dout_10_rsci_dinb_d_reg),
      .dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_10_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_inst_dout_10_rsci_dinb_d_core[63:0]),
      .dout_10_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_inst_dout_10_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_inst
      (
      .dout_11_rsci_dinb_d(dout_11_rsci_dinb_d_reg),
      .dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_11_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_inst_dout_11_rsci_dinb_d_core[63:0]),
      .dout_11_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_inst_dout_11_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_inst
      (
      .dout_12_rsci_dinb_d(dout_12_rsci_dinb_d_reg),
      .dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_12_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_inst_dout_12_rsci_dinb_d_core[63:0]),
      .dout_12_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_inst_dout_12_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_inst
      (
      .dout_13_rsci_dinb_d(dout_13_rsci_dinb_d_reg),
      .dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_13_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_inst_dout_13_rsci_dinb_d_core[63:0]),
      .dout_13_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_inst_dout_13_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_inst
      (
      .dout_14_rsci_dinb_d(dout_14_rsci_dinb_d_reg),
      .dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_14_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_inst_dout_14_rsci_dinb_d_core[63:0]),
      .dout_14_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_inst_dout_14_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_inst
      (
      .dout_15_rsci_dinb_d(dout_15_rsci_dinb_d_reg),
      .dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_15_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_inst_dout_15_rsci_dinb_d_core[63:0]),
      .dout_15_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_inst_dout_15_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_inst
      (
      .dout_16_rsci_dinb_d(dout_16_rsci_dinb_d_reg),
      .dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_16_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_inst_dout_16_rsci_dinb_d_core[63:0]),
      .dout_16_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_inst_dout_16_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_inst
      (
      .dout_17_rsci_dinb_d(dout_17_rsci_dinb_d_reg),
      .dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_17_rsci_dinb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_inst_dout_17_rsci_dinb_d_core[63:0]),
      .dout_17_rsci_iswt0_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_inst_dout_17_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_0_data_rsci_addra_d(tmp_0_data_rsci_addra_d_reg),
      .tmp_0_data_rsci_addrb_d(tmp_0_data_rsci_addrb_d_reg),
      .tmp_0_data_rsci_douta_d(tmp_0_data_rsci_douta_d),
      .tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_0_data_rsci_oswt(reg_tmp_0_data_rsci_oswt_cse),
      .tmp_0_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_addra_d_core[7:0]),
      .tmp_0_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_addrb_d_core[7:0]),
      .tmp_0_data_rsci_douta_d_mxwt(tmp_0_data_rsci_douta_d_mxwt),
      .tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_0_data_rsci_1_inst_tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_0_data_rsci_oswt_pff(WRITE_for_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_1_data_rsci_addra_d(tmp_1_data_rsci_addra_d_reg),
      .tmp_1_data_rsci_addrb_d(tmp_1_data_rsci_addrb_d_reg),
      .tmp_1_data_rsci_douta_d(tmp_1_data_rsci_douta_d),
      .tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_1_data_rsci_oswt(reg_tmp_1_data_rsci_oswt_cse),
      .tmp_1_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_addra_d_core[7:0]),
      .tmp_1_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_addrb_d_core[7:0]),
      .tmp_1_data_rsci_douta_d_mxwt(tmp_1_data_rsci_douta_d_mxwt),
      .tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_1_data_rsci_1_inst_tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_1_data_rsci_oswt_pff(WRITE_for_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_2_data_rsci_addra_d(tmp_2_data_rsci_addra_d_reg),
      .tmp_2_data_rsci_addrb_d(tmp_2_data_rsci_addrb_d_reg),
      .tmp_2_data_rsci_douta_d(tmp_2_data_rsci_douta_d),
      .tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_2_data_rsci_oswt(reg_tmp_2_data_rsci_oswt_cse),
      .tmp_2_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_addra_d_core[7:0]),
      .tmp_2_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_addrb_d_core[7:0]),
      .tmp_2_data_rsci_douta_d_mxwt(tmp_2_data_rsci_douta_d_mxwt),
      .tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_2_data_rsci_1_inst_tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_2_data_rsci_oswt_pff(WRITE_for_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_3_data_rsci_addra_d(tmp_3_data_rsci_addra_d_reg),
      .tmp_3_data_rsci_addrb_d(tmp_3_data_rsci_addrb_d_reg),
      .tmp_3_data_rsci_douta_d(tmp_3_data_rsci_douta_d),
      .tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_3_data_rsci_oswt(reg_tmp_3_data_rsci_oswt_cse),
      .tmp_3_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_addra_d_core[7:0]),
      .tmp_3_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_addrb_d_core[7:0]),
      .tmp_3_data_rsci_douta_d_mxwt(tmp_3_data_rsci_douta_d_mxwt),
      .tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_3_data_rsci_1_inst_tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_3_data_rsci_oswt_pff(WRITE_for_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_4_data_rsci_addra_d(tmp_4_data_rsci_addra_d_reg),
      .tmp_4_data_rsci_addrb_d(tmp_4_data_rsci_addrb_d_reg),
      .tmp_4_data_rsci_douta_d(tmp_4_data_rsci_douta_d),
      .tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_4_data_rsci_oswt(reg_tmp_4_data_rsci_oswt_cse),
      .tmp_4_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_addra_d_core[7:0]),
      .tmp_4_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_addrb_d_core[7:0]),
      .tmp_4_data_rsci_douta_d_mxwt(tmp_4_data_rsci_douta_d_mxwt),
      .tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_4_data_rsci_1_inst_tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_4_data_rsci_oswt_pff(WRITE_for_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_5_data_rsci_addra_d(tmp_5_data_rsci_addra_d_reg),
      .tmp_5_data_rsci_addrb_d(tmp_5_data_rsci_addrb_d_reg),
      .tmp_5_data_rsci_douta_d(tmp_5_data_rsci_douta_d),
      .tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_5_data_rsci_oswt(reg_tmp_5_data_rsci_oswt_cse),
      .tmp_5_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_addra_d_core[7:0]),
      .tmp_5_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_addrb_d_core[7:0]),
      .tmp_5_data_rsci_douta_d_mxwt(tmp_5_data_rsci_douta_d_mxwt),
      .tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_5_data_rsci_1_inst_tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_5_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_6_data_rsci_addra_d(tmp_6_data_rsci_addra_d_reg),
      .tmp_6_data_rsci_addrb_d(tmp_6_data_rsci_addrb_d_reg),
      .tmp_6_data_rsci_douta_d(tmp_6_data_rsci_douta_d),
      .tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_6_data_rsci_oswt(reg_tmp_6_data_rsci_oswt_cse),
      .tmp_6_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_addra_d_core[7:0]),
      .tmp_6_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_addrb_d_core[7:0]),
      .tmp_6_data_rsci_douta_d_mxwt(tmp_6_data_rsci_douta_d_mxwt),
      .tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_6_data_rsci_1_inst_tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_6_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_7_data_rsci_addra_d(tmp_7_data_rsci_addra_d_reg),
      .tmp_7_data_rsci_addrb_d(tmp_7_data_rsci_addrb_d_reg),
      .tmp_7_data_rsci_douta_d(tmp_7_data_rsci_douta_d),
      .tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_7_data_rsci_oswt(reg_tmp_7_data_rsci_oswt_cse),
      .tmp_7_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_addra_d_core[7:0]),
      .tmp_7_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_addrb_d_core[7:0]),
      .tmp_7_data_rsci_douta_d_mxwt(tmp_7_data_rsci_douta_d_mxwt),
      .tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_7_data_rsci_1_inst_tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_7_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_8_data_rsci_addra_d(tmp_8_data_rsci_addra_d_reg),
      .tmp_8_data_rsci_addrb_d(tmp_8_data_rsci_addrb_d_reg),
      .tmp_8_data_rsci_douta_d(tmp_8_data_rsci_douta_d),
      .tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_8_data_rsci_oswt(reg_tmp_8_data_rsci_oswt_cse),
      .tmp_8_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_addra_d_core[7:0]),
      .tmp_8_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_addrb_d_core[7:0]),
      .tmp_8_data_rsci_douta_d_mxwt(tmp_8_data_rsci_douta_d_mxwt),
      .tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_8_data_rsci_1_inst_tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_8_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_9_data_rsci_addra_d(tmp_9_data_rsci_addra_d_reg),
      .tmp_9_data_rsci_addrb_d(tmp_9_data_rsci_addrb_d_reg),
      .tmp_9_data_rsci_douta_d(tmp_9_data_rsci_douta_d),
      .tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_9_data_rsci_oswt(reg_tmp_9_data_rsci_oswt_cse),
      .tmp_9_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_addra_d_core[7:0]),
      .tmp_9_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_addrb_d_core[7:0]),
      .tmp_9_data_rsci_douta_d_mxwt(tmp_9_data_rsci_douta_d_mxwt),
      .tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_9_data_rsci_1_inst_tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_9_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_10_data_rsci_addra_d(tmp_10_data_rsci_addra_d_reg),
      .tmp_10_data_rsci_addrb_d(tmp_10_data_rsci_addrb_d_reg),
      .tmp_10_data_rsci_douta_d(tmp_10_data_rsci_douta_d),
      .tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_10_data_rsci_oswt(reg_tmp_10_data_rsci_oswt_cse),
      .tmp_10_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_addra_d_core[7:0]),
      .tmp_10_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_addrb_d_core[7:0]),
      .tmp_10_data_rsci_douta_d_mxwt(tmp_10_data_rsci_douta_d_mxwt),
      .tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_10_data_rsci_1_inst_tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_10_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_11_data_rsci_addra_d(tmp_11_data_rsci_addra_d_reg),
      .tmp_11_data_rsci_addrb_d(tmp_11_data_rsci_addrb_d_reg),
      .tmp_11_data_rsci_douta_d(tmp_11_data_rsci_douta_d),
      .tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_11_data_rsci_oswt(reg_tmp_11_data_rsci_oswt_cse),
      .tmp_11_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_addra_d_core[7:0]),
      .tmp_11_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_addrb_d_core[7:0]),
      .tmp_11_data_rsci_douta_d_mxwt(tmp_11_data_rsci_douta_d_mxwt),
      .tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_11_data_rsci_1_inst_tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_11_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_12_data_rsci_addra_d(tmp_12_data_rsci_addra_d_reg),
      .tmp_12_data_rsci_addrb_d(tmp_12_data_rsci_addrb_d_reg),
      .tmp_12_data_rsci_douta_d(tmp_12_data_rsci_douta_d),
      .tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_12_data_rsci_oswt(reg_tmp_12_data_rsci_oswt_cse),
      .tmp_12_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_addra_d_core[7:0]),
      .tmp_12_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_addrb_d_core[7:0]),
      .tmp_12_data_rsci_douta_d_mxwt(tmp_12_data_rsci_douta_d_mxwt),
      .tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_12_data_rsci_1_inst_tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_12_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_13_data_rsci_addra_d(tmp_13_data_rsci_addra_d_reg),
      .tmp_13_data_rsci_addrb_d(tmp_13_data_rsci_addrb_d_reg),
      .tmp_13_data_rsci_douta_d(tmp_13_data_rsci_douta_d),
      .tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_13_data_rsci_oswt(reg_tmp_13_data_rsci_oswt_cse),
      .tmp_13_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_addra_d_core[7:0]),
      .tmp_13_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_addrb_d_core[7:0]),
      .tmp_13_data_rsci_douta_d_mxwt(tmp_13_data_rsci_douta_d_mxwt),
      .tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_13_data_rsci_1_inst_tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_13_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_14_data_rsci_addra_d(tmp_14_data_rsci_addra_d_reg),
      .tmp_14_data_rsci_addrb_d(tmp_14_data_rsci_addrb_d_reg),
      .tmp_14_data_rsci_douta_d(tmp_14_data_rsci_douta_d),
      .tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_14_data_rsci_oswt(reg_tmp_14_data_rsci_oswt_cse),
      .tmp_14_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_addra_d_core[7:0]),
      .tmp_14_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_addrb_d_core[7:0]),
      .tmp_14_data_rsci_douta_d_mxwt(tmp_14_data_rsci_douta_d_mxwt),
      .tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_14_data_rsci_1_inst_tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_14_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_15_data_rsci_addra_d(tmp_15_data_rsci_addra_d_reg),
      .tmp_15_data_rsci_addrb_d(tmp_15_data_rsci_addrb_d_reg),
      .tmp_15_data_rsci_douta_d(tmp_15_data_rsci_douta_d),
      .tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_15_data_rsci_oswt(reg_tmp_15_data_rsci_oswt_cse),
      .tmp_15_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_addra_d_core[7:0]),
      .tmp_15_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_addrb_d_core[7:0]),
      .tmp_15_data_rsci_douta_d_mxwt(tmp_15_data_rsci_douta_d_mxwt),
      .tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_15_data_rsci_1_inst_tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_15_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_16_data_rsci_addra_d(tmp_16_data_rsci_addra_d_reg),
      .tmp_16_data_rsci_addrb_d(tmp_16_data_rsci_addrb_d_reg),
      .tmp_16_data_rsci_douta_d(tmp_16_data_rsci_douta_d),
      .tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_16_data_rsci_oswt(reg_tmp_16_data_rsci_oswt_cse),
      .tmp_16_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_addra_d_core[7:0]),
      .tmp_16_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_addrb_d_core[7:0]),
      .tmp_16_data_rsci_douta_d_mxwt(tmp_16_data_rsci_douta_d_mxwt),
      .tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_16_data_rsci_1_inst_tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_16_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .tmp_17_data_rsci_addra_d(tmp_17_data_rsci_addra_d_reg),
      .tmp_17_data_rsci_addrb_d(tmp_17_data_rsci_addrb_d_reg),
      .tmp_17_data_rsci_douta_d(tmp_17_data_rsci_douta_d),
      .tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .tmp_17_data_rsci_oswt(reg_tmp_17_data_rsci_oswt_cse),
      .tmp_17_data_rsci_addra_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_addra_d_core[7:0]),
      .tmp_17_data_rsci_addrb_d_core(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_addrb_d_core[7:0]),
      .tmp_17_data_rsci_douta_d_mxwt(tmp_17_data_rsci_douta_d_mxwt),
      .tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct[0:0]),
      .tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct(nl_WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_tmp_17_data_rsci_1_inst_tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_core_psct[0:0]),
      .tmp_17_data_rsci_oswt_pff(WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_rls_obj_inst
      (
      .dout_17_rsc_rls_lz(dout_17_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_17_rsc_rls_obj_iswt0(reg_dout_17_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_17_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_17_rsc_req_vz(dout_17_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_17_rsc_req_obj_oswt(reg_dout_17_rsc_req_obj_oswt_cse),
      .dout_17_rsc_req_obj_wen_comp(dout_17_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_rls_obj_inst
      (
      .dout_16_rsc_rls_lz(dout_16_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_16_rsc_rls_obj_iswt0(reg_dout_16_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_16_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_16_rsc_req_vz(dout_16_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_16_rsc_req_obj_oswt(reg_dout_16_rsc_req_obj_oswt_cse),
      .dout_16_rsc_req_obj_wen_comp(dout_16_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_rls_obj_inst
      (
      .dout_15_rsc_rls_lz(dout_15_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_15_rsc_rls_obj_iswt0(reg_dout_15_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_15_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_15_rsc_req_vz(dout_15_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_15_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_15_rsc_req_obj_wen_comp(dout_15_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_rls_obj_inst
      (
      .dout_14_rsc_rls_lz(dout_14_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_14_rsc_rls_obj_iswt0(reg_dout_14_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_14_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_14_rsc_req_vz(dout_14_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_14_rsc_req_obj_oswt(reg_dout_14_rsc_req_obj_oswt_cse),
      .dout_14_rsc_req_obj_wen_comp(dout_14_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_rls_obj_inst
      (
      .dout_13_rsc_rls_lz(dout_13_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_13_rsc_rls_obj_iswt0(reg_dout_13_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_13_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_13_rsc_req_vz(dout_13_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_13_rsc_req_obj_oswt(reg_dout_13_rsc_req_obj_oswt_cse),
      .dout_13_rsc_req_obj_wen_comp(dout_13_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_rls_obj_inst
      (
      .dout_12_rsc_rls_lz(dout_12_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_12_rsc_rls_obj_iswt0(reg_dout_12_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_12_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_12_rsc_req_vz(dout_12_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_12_rsc_req_obj_oswt(reg_dout_12_rsc_req_obj_oswt_cse),
      .dout_12_rsc_req_obj_wen_comp(dout_12_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_rls_obj_inst
      (
      .dout_11_rsc_rls_lz(dout_11_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_11_rsc_rls_obj_iswt0(reg_dout_11_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_11_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_11_rsc_req_vz(dout_11_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_11_rsc_req_obj_oswt(reg_dout_11_rsc_req_obj_oswt_cse),
      .dout_11_rsc_req_obj_wen_comp(dout_11_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_rls_obj_inst
      (
      .dout_10_rsc_rls_lz(dout_10_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_10_rsc_rls_obj_iswt0(reg_dout_10_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_10_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_10_rsc_req_vz(dout_10_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_10_rsc_req_obj_oswt(reg_dout_10_rsc_req_obj_oswt_cse),
      .dout_10_rsc_req_obj_wen_comp(dout_10_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_rls_obj_inst
      (
      .dout_9_rsc_rls_lz(dout_9_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_9_rsc_rls_obj_iswt0(reg_dout_9_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_9_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_9_rsc_req_vz(dout_9_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_9_rsc_req_obj_oswt(reg_dout_9_rsc_req_obj_oswt_cse),
      .dout_9_rsc_req_obj_wen_comp(dout_9_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_rls_obj_inst
      (
      .dout_8_rsc_rls_lz(dout_8_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_8_rsc_rls_obj_iswt0(reg_dout_8_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_8_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_8_rsc_req_vz(dout_8_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_8_rsc_req_obj_oswt(reg_dout_8_rsc_req_obj_oswt_cse),
      .dout_8_rsc_req_obj_wen_comp(dout_8_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_rls_obj_inst
      (
      .dout_7_rsc_rls_lz(dout_7_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_7_rsc_rls_obj_iswt0(reg_dout_7_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_7_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_7_rsc_req_vz(dout_7_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_7_rsc_req_obj_oswt(reg_dout_7_rsc_req_obj_oswt_cse),
      .dout_7_rsc_req_obj_wen_comp(dout_7_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_rls_obj_inst
      (
      .dout_6_rsc_rls_lz(dout_6_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_6_rsc_rls_obj_iswt0(reg_dout_6_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_6_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_6_rsc_req_vz(dout_6_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_6_rsc_req_obj_oswt(reg_dout_6_rsc_req_obj_oswt_cse),
      .dout_6_rsc_req_obj_wen_comp(dout_6_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_rls_obj_inst
      (
      .dout_5_rsc_rls_lz(dout_5_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_5_rsc_rls_obj_iswt0(reg_dout_5_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_5_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_5_rsc_req_vz(dout_5_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_5_rsc_req_obj_oswt(reg_dout_5_rsc_req_obj_oswt_cse),
      .dout_5_rsc_req_obj_wen_comp(dout_5_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_rls_obj_inst
      (
      .dout_4_rsc_rls_lz(dout_4_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_4_rsc_rls_obj_iswt0(reg_dout_4_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_4_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_4_rsc_req_vz(dout_4_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_4_rsc_req_obj_oswt(reg_dout_4_rsc_req_obj_oswt_cse),
      .dout_4_rsc_req_obj_wen_comp(dout_4_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_rls_obj_inst
      (
      .dout_3_rsc_rls_lz(dout_3_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_3_rsc_rls_obj_iswt0(reg_dout_3_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_3_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_3_rsc_req_vz(dout_3_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_3_rsc_req_obj_oswt(reg_dout_3_rsc_req_obj_oswt_cse),
      .dout_3_rsc_req_obj_wen_comp(dout_3_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_rls_obj_inst
      (
      .dout_2_rsc_rls_lz(dout_2_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_2_rsc_rls_obj_iswt0(reg_dout_2_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_2_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_2_rsc_req_vz(dout_2_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_2_rsc_req_obj_oswt(reg_dout_2_rsc_req_obj_oswt_cse),
      .dout_2_rsc_req_obj_wen_comp(dout_2_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_rls_obj_inst
      (
      .dout_1_rsc_rls_lz(dout_1_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_1_rsc_rls_obj_iswt0(reg_dout_1_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_1_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_1_rsc_req_vz(dout_1_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_1_rsc_req_obj_oswt(reg_dout_1_rsc_req_obj_oswt_cse),
      .dout_1_rsc_req_obj_wen_comp(dout_1_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_rls_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_rls_obj_inst
      (
      .dout_0_rsc_rls_lz(dout_0_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_0_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_iswt0_cse)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_dout_0_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_0_rsc_req_vz(dout_0_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_0_rsc_req_obj_oswt(reg_dout_0_rsc_req_obj_oswt_cse),
      .dout_0_rsc_req_obj_wen_comp(dout_0_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_staller WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .core_wten(core_wten),
      .dout_17_rsc_req_obj_wen_comp(dout_17_rsc_req_obj_wen_comp),
      .dout_16_rsc_req_obj_wen_comp(dout_16_rsc_req_obj_wen_comp),
      .dout_15_rsc_req_obj_wen_comp(dout_15_rsc_req_obj_wen_comp),
      .dout_14_rsc_req_obj_wen_comp(dout_14_rsc_req_obj_wen_comp),
      .dout_13_rsc_req_obj_wen_comp(dout_13_rsc_req_obj_wen_comp),
      .dout_12_rsc_req_obj_wen_comp(dout_12_rsc_req_obj_wen_comp),
      .dout_11_rsc_req_obj_wen_comp(dout_11_rsc_req_obj_wen_comp),
      .dout_10_rsc_req_obj_wen_comp(dout_10_rsc_req_obj_wen_comp),
      .dout_9_rsc_req_obj_wen_comp(dout_9_rsc_req_obj_wen_comp),
      .dout_8_rsc_req_obj_wen_comp(dout_8_rsc_req_obj_wen_comp),
      .dout_7_rsc_req_obj_wen_comp(dout_7_rsc_req_obj_wen_comp),
      .dout_6_rsc_req_obj_wen_comp(dout_6_rsc_req_obj_wen_comp),
      .dout_5_rsc_req_obj_wen_comp(dout_5_rsc_req_obj_wen_comp),
      .dout_4_rsc_req_obj_wen_comp(dout_4_rsc_req_obj_wen_comp),
      .dout_3_rsc_req_obj_wen_comp(dout_3_rsc_req_obj_wen_comp),
      .dout_2_rsc_req_obj_wen_comp(dout_2_rsc_req_obj_wen_comp),
      .dout_1_rsc_req_obj_wen_comp(dout_1_rsc_req_obj_wen_comp),
      .dout_0_rsc_req_obj_wen_comp(dout_0_rsc_req_obj_wen_comp)
    );
  assign and_206_cse = core_wen & main_stage_0_2 & equal_tmp_50;
  assign and_208_cse = core_wen & main_stage_0_2 & equal_tmp_48;
  assign and_210_cse = core_wen & main_stage_0_2 & equal_tmp_46;
  assign and_212_cse = core_wen & main_stage_0_2 & equal_tmp_44;
  assign and_214_cse = core_wen & main_stage_0_2 & equal_tmp_42;
  assign and_216_cse = core_wen & main_stage_0_2 & equal_tmp_40;
  assign and_218_cse = core_wen & main_stage_0_2 & equal_tmp_38;
  assign and_220_cse = core_wen & main_stage_0_2 & equal_tmp_36;
  assign and_222_cse = core_wen & main_stage_0_2 & equal_tmp_34;
  assign and_224_cse = core_wen & main_stage_0_2 & equal_tmp_32;
  assign and_226_cse = core_wen & main_stage_0_2 & equal_tmp_30;
  assign and_228_cse = core_wen & main_stage_0_2 & equal_tmp_28;
  assign and_230_cse = core_wen & main_stage_0_2 & equal_tmp_26;
  assign and_232_cse = core_wen & main_stage_0_2 & equal_tmp_24;
  assign and_234_cse = core_wen & main_stage_0_2 & equal_tmp_22;
  assign and_236_cse = core_wen & main_stage_0_2 & equal_tmp_20;
  assign and_238_cse = core_wen & main_stage_0_2 & equal_tmp_18;
  assign or_358_nl = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1:0]!=2'b10);
  assign or_359_nl = (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]);
  assign mux_149_nl = MUX_s_1_2_2((or_359_nl), (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]),
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign mux_150_nl = MUX_s_1_2_2((mux_149_nl), (or_358_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_if_nor_rmff = ~((mux_150_nl) | or_dcpl_246);
  assign WRITE_x_idx_mux_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_0_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign and_168_nl = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1:0]==2'b11);
  assign nor_116_nl = ~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0])) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]));
  assign mux_151_nl = MUX_s_1_2_2((nor_116_nl), (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]),
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign mux_152_nl = MUX_s_1_2_2((mux_151_nl), (and_168_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_if_nor_rmff = ~((~ (mux_152_nl)) | or_dcpl_246);
  assign WRITE_x_idx_mux_1_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_1_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign or_375_nl = (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2])
      | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3])
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]);
  assign mux_153_nl = MUX_s_1_2_2(or_tmp_75, (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]),
      WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]);
  assign mux_154_nl = MUX_s_1_2_2((~ (mux_153_nl)), (or_375_nl), lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]);
  assign mux_155_nl = MUX_s_1_2_2((mux_154_nl), or_dcpl_213, WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_if_nor_rmff = ~((mux_155_nl) | or_dcpl_260);
  assign WRITE_x_idx_mux_2_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_2_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign mux_156_nl = MUX_s_1_2_2((lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]),
      or_tmp_75, WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]);
  assign nor_114_nl = ~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0])) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2])
      | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3])
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]));
  assign mux_157_nl = MUX_s_1_2_2((nor_114_nl), (mux_156_nl), lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]);
  assign mux_158_nl = MUX_s_1_2_2((mux_157_nl), nor_tmp_21, WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_if_nor_rmff = ~((~ (mux_158_nl)) | or_dcpl_260);
  assign WRITE_x_idx_mux_3_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_3_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign or_388_nl = (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2])
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3])
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]);
  assign mux_159_nl = MUX_s_1_2_2((or_388_nl), or_dcpl_213, lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign mux_160_nl = MUX_s_1_2_2(or_dcpl_214, (mux_159_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_if_nor_rmff = ~((mux_160_nl) | or_dcpl_232);
  assign WRITE_x_idx_mux_4_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_4_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign nor_113_nl = ~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0])) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2])
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3])
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]));
  assign mux_161_nl = MUX_s_1_2_2((nor_113_nl), nor_tmp_21, lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign and_166_nl = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2:0]==3'b111);
  assign mux_162_nl = MUX_s_1_2_2((and_166_nl), (mux_161_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_if_nor_rmff = ~((~ (mux_162_nl)) | or_dcpl_232);
  assign WRITE_x_idx_mux_5_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_5_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign or_400_nl = (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]))
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]);
  assign nor_111_nl = ~((~((WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]))
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])))
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]));
  assign mux_163_nl = MUX_s_1_2_2((nor_111_nl), (or_400_nl), lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]);
  assign mux_164_nl = MUX_s_1_2_2(or_tmp_82, (mux_163_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_else_if_nor_rmff = ~((mux_164_nl) | or_dcpl_279);
  assign WRITE_x_idx_mux_6_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_6_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]);
  assign or_408_nl = (~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0])) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]))
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])))
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]);
  assign nor_110_nl = ~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0])) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]))
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]));
  assign mux_165_nl = MUX_s_1_2_2((nor_110_nl), (or_408_nl), lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]);
  assign mux_166_nl = MUX_s_1_2_2(nor_tmp_23, (mux_165_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_else_else_if_nor_rmff = ~((~ (mux_166_nl))
      | or_dcpl_279);
  assign WRITE_x_idx_mux_7_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_7_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]);
  assign or_415_nl = (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1])) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0])
      | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]));
  assign or_416_nl = (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])
      | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3])) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]);
  assign mux_167_nl = MUX_s_1_2_2((or_416_nl), or_tmp_82, lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign mux_168_nl = MUX_s_1_2_2((mux_167_nl), (or_415_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_else_else_else_if_nor_rmff = ~((mux_168_nl)
      | or_dcpl_286);
  assign WRITE_x_idx_mux_8_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_8_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign and_164_nl = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]) & (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0])
      & (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]);
  assign nor_108_nl = ~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0])) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])
      | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3])) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]));
  assign mux_169_nl = MUX_s_1_2_2((nor_108_nl), nor_tmp_23, lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign mux_170_nl = MUX_s_1_2_2((mux_169_nl), (and_164_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_else_else_else_else_if_nor_rmff = ~((~
      (mux_170_nl)) | or_dcpl_286);
  assign WRITE_x_idx_mux_9_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_9_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign or_426_nl = (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2])
      | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]))
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]);
  assign mux_172_nl = MUX_s_1_2_2(mux_tmp_42, nor_tmp_25, WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]);
  assign mux_173_nl = MUX_s_1_2_2((~ (mux_172_nl)), (or_426_nl), lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]);
  assign mux_174_nl = MUX_s_1_2_2((mux_173_nl), or_tmp_90, WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_else_else_else_else_else_if_nor_rmff
      = ~((mux_174_nl) | or_dcpl_293);
  assign WRITE_x_idx_mux_10_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_10_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign mux_175_nl = MUX_s_1_2_2(nor_tmp_25, mux_tmp_42, WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]);
  assign nor_107_nl = ~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0])) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2])
      | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]))
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]));
  assign mux_176_nl = MUX_s_1_2_2((nor_107_nl), (mux_175_nl), lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]);
  assign mux_177_nl = MUX_s_1_2_2((mux_176_nl), nor_tmp_26, WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff
      = ~((~ (mux_177_nl)) | or_dcpl_293);
  assign WRITE_x_idx_mux_11_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_11_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign or_433_nl = (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2])
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]))
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]);
  assign mux_178_nl = MUX_s_1_2_2((or_433_nl), or_tmp_90, lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign or_435_nl = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1:0]!=2'b10) |
      (~ nor_tmp_25);
  assign mux_179_nl = MUX_s_1_2_2((or_435_nl), (mux_178_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff
      = ~((mux_179_nl) | or_dcpl_278);
  assign WRITE_x_idx_mux_12_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_12_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign nor_106_nl = ~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0])) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2])
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]))
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]));
  assign mux_180_nl = MUX_s_1_2_2((nor_106_nl), nor_tmp_26, lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign and_161_nl = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3:0]==4'b1111);
  assign mux_181_nl = MUX_s_1_2_2((and_161_nl), (mux_180_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff
      = ~((~ (mux_181_nl)) | or_dcpl_278);
  assign WRITE_x_idx_mux_13_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_13_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign or_442_nl = (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]))
      | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3])) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]);
  assign nor_104_nl = ~((~((WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]))
      | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3])) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])))
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]));
  assign mux_182_nl = MUX_s_1_2_2((nor_104_nl), (or_442_nl), lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]);
  assign mux_183_nl = MUX_s_1_2_2(or_tmp_101, (mux_182_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff
      = ~((mux_183_nl) | or_dcpl_302);
  assign WRITE_x_idx_mux_14_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_14_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]);
  assign or_449_nl = ((WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]) & (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])
      & (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]) & (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])))
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]);
  assign nor_103_nl = ~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0])) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]))
      | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3])) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]));
  assign mux_184_nl = MUX_s_1_2_2((nor_103_nl), (or_449_nl), lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]);
  assign mux_185_nl = MUX_s_1_2_2(nor_tmp_28, (mux_184_nl), WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff
      = ~((~ (mux_185_nl)) | or_dcpl_302);
  assign WRITE_x_idx_mux_15_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_15_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]);
  assign or_454_nl = WRITE_for_y_idx_slc_WRITE_for_y_idx_4_0_0_itm_3 | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]))
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]);
  assign mux_186_nl = MUX_s_1_2_2((or_454_nl), or_tmp_101, lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff
      = ~((mux_186_nl) | or_dcpl_307);
  assign WRITE_x_idx_mux_16_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, io_write_dout_16_copy_ndx_6_0_lpi_1_mx0,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign nor_102_nl = ~((~ WRITE_for_y_idx_slc_WRITE_for_y_idx_4_0_0_itm_3) | (~
      (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]));
  assign mux_187_nl = MUX_s_1_2_2((nor_102_nl), nor_tmp_28, lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff
      = ~((~ (mux_187_nl)) | or_dcpl_307);
  assign WRITE_x_idx_mux_17_rmff = MUX_v_7_2_2(WRITE_x_idx_6_0_lpi_1_dfm_5, mux_53_tmp,
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign mux_130_cse = MUX_s_1_2_2((~ exit_WRITE_lpi_1_dfm_4), lfst_exit_WRITE_lpi_1,
      or_2_tmp_1);
  assign or_3_tmp = equal_tmp_73 | equal_tmp_74 | equal_tmp_75 | equal_tmp_76 | equal_tmp_77
      | equal_tmp_78 | equal_tmp_79 | equal_tmp_80 | equal_tmp_81 | equal_tmp_82
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_3_tmp = MUX1HOT_v_7_3_2(io_write_dout_0_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_0_copy_ndx_6_0_sva_4, io_write_dout_0_copy_ndx_6_0_lpi_1, {nor_dfs_3
      , equal_tmp_72 , or_3_tmp});
  assign io_write_dout_0_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_0_copy_ndx_6_0_lpi_1,
      mux1h_3_tmp, main_stage_0_3);
  assign or_4_tmp = nor_dfs_3 | equal_tmp_74 | equal_tmp_75 | equal_tmp_76 | equal_tmp_77
      | equal_tmp_78 | equal_tmp_79 | equal_tmp_80 | equal_tmp_81 | equal_tmp_82
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_4_tmp = MUX1HOT_v_7_3_2(io_write_dout_1_copy_ndx_6_0_lpi_1, io_write_dout_1_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_1_copy_ndx_6_0_sva_4, {or_4_tmp , equal_tmp_72 , equal_tmp_73});
  assign io_write_dout_1_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_1_copy_ndx_6_0_lpi_1,
      mux1h_4_tmp, main_stage_0_3);
  assign or_5_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_75 | equal_tmp_76 | equal_tmp_77
      | equal_tmp_78 | equal_tmp_79 | equal_tmp_80 | equal_tmp_81 | equal_tmp_82
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_5_tmp = MUX1HOT_v_7_3_2(io_write_dout_2_copy_ndx_6_0_lpi_1, io_write_dout_2_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_2_copy_ndx_6_0_sva_4, {or_5_tmp , equal_tmp_73 , equal_tmp_74});
  assign io_write_dout_2_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_2_copy_ndx_6_0_lpi_1,
      mux1h_5_tmp, main_stage_0_3);
  assign or_6_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_76 | equal_tmp_77
      | equal_tmp_78 | equal_tmp_79 | equal_tmp_80 | equal_tmp_81 | equal_tmp_82
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_6_tmp = MUX1HOT_v_7_3_2(io_write_dout_3_copy_ndx_6_0_lpi_1, io_write_dout_3_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_3_copy_ndx_6_0_sva_4, {or_6_tmp , equal_tmp_74 , equal_tmp_75});
  assign io_write_dout_3_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_3_copy_ndx_6_0_lpi_1,
      mux1h_6_tmp, main_stage_0_3);
  assign or_7_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_77
      | equal_tmp_78 | equal_tmp_79 | equal_tmp_80 | equal_tmp_81 | equal_tmp_82
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_7_tmp = MUX1HOT_v_7_3_2(io_write_dout_4_copy_ndx_6_0_lpi_1, io_write_dout_4_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_4_copy_ndx_6_0_sva_4, {or_7_tmp , equal_tmp_75 , equal_tmp_76});
  assign io_write_dout_4_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_4_copy_ndx_6_0_lpi_1,
      mux1h_7_tmp, main_stage_0_3);
  assign or_8_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_78 | equal_tmp_79 | equal_tmp_80 | equal_tmp_81 | equal_tmp_82
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_8_tmp = MUX1HOT_v_7_3_2(io_write_dout_5_copy_ndx_6_0_lpi_1, io_write_dout_5_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_5_copy_ndx_6_0_sva_4, {or_8_tmp , equal_tmp_76 , equal_tmp_77});
  assign io_write_dout_5_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_5_copy_ndx_6_0_lpi_1,
      mux1h_8_tmp, main_stage_0_3);
  assign or_9_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_79 | equal_tmp_80 | equal_tmp_81 | equal_tmp_82
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_9_tmp = MUX1HOT_v_7_3_2(io_write_dout_6_copy_ndx_6_0_lpi_1, io_write_dout_6_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_6_copy_ndx_6_0_sva_4, {or_9_tmp , equal_tmp_77 , equal_tmp_78});
  assign io_write_dout_6_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_6_copy_ndx_6_0_lpi_1,
      mux1h_9_tmp, main_stage_0_3);
  assign or_10_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_80 | equal_tmp_81 | equal_tmp_82
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_10_tmp = MUX1HOT_v_7_3_2(io_write_dout_7_copy_ndx_6_0_lpi_1, io_write_dout_7_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_7_copy_ndx_6_0_sva_4, {or_10_tmp , equal_tmp_78 , equal_tmp_79});
  assign io_write_dout_7_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_7_copy_ndx_6_0_lpi_1,
      mux1h_10_tmp, main_stage_0_3);
  assign or_11_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_78 | equal_tmp_81 | equal_tmp_82
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_11_tmp = MUX1HOT_v_7_3_2(io_write_dout_8_copy_ndx_6_0_lpi_1, io_write_dout_8_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_8_copy_ndx_6_0_sva_4, {or_11_tmp , equal_tmp_79 , equal_tmp_80});
  assign io_write_dout_8_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_8_copy_ndx_6_0_lpi_1,
      mux1h_11_tmp, main_stage_0_3);
  assign or_12_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_78 | equal_tmp_79 | equal_tmp_82
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_12_tmp = MUX1HOT_v_7_3_2(io_write_dout_9_copy_ndx_6_0_lpi_1, io_write_dout_9_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_9_copy_ndx_6_0_sva_4, {or_12_tmp , equal_tmp_80 , equal_tmp_81});
  assign io_write_dout_9_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_9_copy_ndx_6_0_lpi_1,
      mux1h_12_tmp, main_stage_0_3);
  assign or_13_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_78 | equal_tmp_79 | equal_tmp_80
      | equal_tmp_83 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_13_tmp = MUX1HOT_v_7_3_2(io_write_dout_10_copy_ndx_6_0_lpi_1, io_write_dout_10_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_10_copy_ndx_6_0_sva_4, {or_13_tmp , equal_tmp_81 , equal_tmp_82});
  assign io_write_dout_10_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_10_copy_ndx_6_0_lpi_1,
      mux1h_13_tmp, main_stage_0_3);
  assign or_14_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_78 | equal_tmp_79 | equal_tmp_80
      | equal_tmp_81 | equal_tmp_84 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_14_tmp = MUX1HOT_v_7_3_2(io_write_dout_11_copy_ndx_6_0_lpi_1, io_write_dout_11_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_11_copy_ndx_6_0_sva_4, {or_14_tmp , equal_tmp_82 , equal_tmp_83});
  assign io_write_dout_11_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_11_copy_ndx_6_0_lpi_1,
      mux1h_14_tmp, main_stage_0_3);
  assign or_15_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_78 | equal_tmp_79 | equal_tmp_80
      | equal_tmp_81 | equal_tmp_82 | equal_tmp_85 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_15_tmp = MUX1HOT_v_7_3_2(io_write_dout_12_copy_ndx_6_0_lpi_1, io_write_dout_12_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_12_copy_ndx_6_0_sva_4, {or_15_tmp , equal_tmp_83 , equal_tmp_84});
  assign io_write_dout_12_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_12_copy_ndx_6_0_lpi_1,
      mux1h_15_tmp, main_stage_0_3);
  assign or_16_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_78 | equal_tmp_79 | equal_tmp_80
      | equal_tmp_81 | equal_tmp_82 | equal_tmp_83 | equal_tmp_86 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_16_tmp = MUX1HOT_v_7_3_2(io_write_dout_13_copy_ndx_6_0_lpi_1, io_write_dout_13_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_13_copy_ndx_6_0_sva_4, {or_16_tmp , equal_tmp_84 , equal_tmp_85});
  assign io_write_dout_13_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_13_copy_ndx_6_0_lpi_1,
      mux1h_16_tmp, main_stage_0_3);
  assign or_17_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_78 | equal_tmp_79 | equal_tmp_80
      | equal_tmp_81 | equal_tmp_82 | equal_tmp_83 | equal_tmp_84 | equal_tmp_87
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_17_tmp = MUX1HOT_v_7_3_2(io_write_dout_14_copy_ndx_6_0_lpi_1, io_write_dout_14_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_14_copy_ndx_6_0_sva_4, {or_17_tmp , equal_tmp_85 , equal_tmp_86});
  assign io_write_dout_14_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_14_copy_ndx_6_0_lpi_1,
      mux1h_17_tmp, main_stage_0_3);
  assign or_18_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_78 | equal_tmp_79 | equal_tmp_80
      | equal_tmp_81 | equal_tmp_82 | equal_tmp_83 | equal_tmp_84 | equal_tmp_85
      | equal_tmp_88 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_18_tmp = MUX1HOT_v_7_3_2(io_write_dout_15_copy_ndx_6_0_lpi_1, io_write_dout_15_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_15_copy_ndx_6_0_sva_4, {or_18_tmp , equal_tmp_86 , equal_tmp_87});
  assign io_write_dout_15_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_15_copy_ndx_6_0_lpi_1,
      mux1h_18_tmp, main_stage_0_3);
  assign or_19_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_78 | equal_tmp_79 | equal_tmp_80
      | equal_tmp_81 | equal_tmp_82 | equal_tmp_83 | equal_tmp_84 | equal_tmp_85
      | equal_tmp_86 | equal_tmp_89 | nor_tmp_30;
  assign mux1h_19_tmp = MUX1HOT_v_7_3_2(io_write_dout_16_copy_ndx_6_0_lpi_1, io_write_dout_16_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_16_copy_ndx_6_0_sva_4, {or_19_tmp , equal_tmp_87 , equal_tmp_88});
  assign io_write_dout_16_copy_ndx_6_0_lpi_1_mx0 = MUX_v_7_2_2(io_write_dout_16_copy_ndx_6_0_lpi_1,
      mux1h_19_tmp, main_stage_0_3);
  assign or_20_tmp = nor_dfs_3 | equal_tmp_72 | equal_tmp_73 | equal_tmp_74 | equal_tmp_75
      | equal_tmp_76 | equal_tmp_77 | equal_tmp_78 | equal_tmp_79 | equal_tmp_80
      | equal_tmp_81 | equal_tmp_82 | equal_tmp_83 | equal_tmp_84 | equal_tmp_85
      | equal_tmp_86 | equal_tmp_87 | nor_tmp_30;
  assign or_568_nl = (~ main_stage_0_3) | or_20_tmp;
  assign and_190_nl = equal_tmp_88 & main_stage_0_3;
  assign and_191_nl = equal_tmp_89 & main_stage_0_3;
  assign mux_53_tmp = MUX1HOT_v_7_3_2(io_write_dout_17_copy_ndx_6_0_lpi_1, io_write_dout_17_copy_ndx_6_0_lpi_1_dfm_4,
      io_write_dout_17_copy_ndx_6_0_sva_4, {(or_568_nl) , (and_190_nl) , (and_191_nl)});
  assign and_169_nl = ((mux1h_78_tmp!=5'b00000)) & main_stage_0_2;
  assign lfst_exit_io_write_dout_17_copy_lpi_1_dfm = MUX_v_5_2_2(5'b00000, mux1h_78_tmp,
      (and_169_nl));
  assign nor_19_tmp = ~(equal_tmp_18 | equal_tmp_20 | equal_tmp_22 | equal_tmp_24
      | equal_tmp_26 | equal_tmp_28 | equal_tmp_30 | equal_tmp_32 | equal_tmp_34
      | equal_tmp_36 | equal_tmp_38 | equal_tmp_40 | equal_tmp_42 | equal_tmp_44
      | equal_tmp_46 | equal_tmp_48 | equal_tmp_50 | equal_tmp_52 | nor_tmp_1);
  assign nl_WRITE_for_acc_nl = conv_u2s_4_5(WRITE_for_y_idx_4_0_sva_1[4:1]) + 5'b10111;
  assign WRITE_for_acc_nl = nl_WRITE_for_acc_nl[4:0];
  assign WRITE_for_acc_itm_4_1 = readslicef_5_1_4((WRITE_for_acc_nl));
  assign nl_WRITE_for_y_idx_4_0_sva_1 = WRITE_for_y_idx_4_0_lpi_1_dfm + 5'b1;
  assign WRITE_for_y_idx_4_0_sva_1 = nl_WRITE_for_y_idx_4_0_sva_1[4:0];
  assign for_for_and_1_nl = lfst_exit_WRITE_lpi_1_mx0 & for_unequal_tmp;
  assign WRITE_for_y_idx_4_0_lpi_1_dfm = MUX_v_5_2_2(5'b00000, mux1h_77_tmp, (for_for_and_1_nl));
  assign nor_tmp_31 = ~((~(WRITE_for_slc_WRITE_for_acc_4_svs_2 | exit_WRITE_sva_2))
      | or_2_tmp_1);
  assign nor_257_nl = ~(or_2_tmp_1 | nor_tmp_31);
  assign mux1h_77_tmp = MUX1HOT_v_5_3_2(({{4{exit_WRITE_sva_2}}, exit_WRITE_sva_2}),
      WRITE_for_y_idx_4_0_lpi_3, WRITE_for_y_idx_4_0_sva_6, {(nor_257_nl) , or_2_tmp_1
      , nor_tmp_31});
  assign or_472_nl = (~ main_stage_0_2) | or_2_tmp_1;
  assign lfst_exit_WRITE_lpi_1_mx0 = MUX_s_1_2_2((~ exit_WRITE_lpi_1_dfm_4), lfst_exit_WRITE_lpi_1,
      or_472_nl);
  assign for_unequal_tmp = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm!=5'b00000);
  assign or_732_tmp = (((mux_53_tmp!=7'b1000001)) & equal_tmp_52) | (unequal_tmp
      & equal_tmp_18) | (unequal_tmp_1 & equal_tmp_20) | (unequal_tmp_2 & equal_tmp_22)
      | (unequal_tmp_3 & equal_tmp_24) | (unequal_tmp_4 & equal_tmp_26) | (unequal_tmp_5
      & equal_tmp_28) | (unequal_tmp_6 & equal_tmp_30) | (unequal_tmp_7 & equal_tmp_32)
      | (unequal_tmp_8 & equal_tmp_34) | (unequal_tmp_9 & equal_tmp_36) | (unequal_tmp_10
      & equal_tmp_38) | (unequal_tmp_11 & equal_tmp_40) | (unequal_tmp_12 & equal_tmp_42)
      | (unequal_tmp_13 & equal_tmp_44) | (unequal_tmp_14 & equal_tmp_46) | (unequal_tmp_15
      & equal_tmp_48) | (unequal_tmp_16 & equal_tmp_50) | nor_tmp_1;
  assign for_mux_3_nl = MUX_v_2_2_2(2'b1, 2'b10, exit_WRITE_lpi_1_dfm_4);
  assign nand_17_nl = ~((mux_53_tmp==7'b1000001));
  assign and_202_nl = nor_19_tmp & (~ or_732_tmp);
  assign and_79_nl = (~ unequal_tmp) & equal_tmp_18 & (~ or_732_tmp);
  assign and_81_nl = (~ unequal_tmp_1) & equal_tmp_20 & (~ or_732_tmp);
  assign and_83_nl = (~ unequal_tmp_2) & equal_tmp_22 & (~ or_732_tmp);
  assign and_85_nl = (~ unequal_tmp_3) & equal_tmp_24 & (~ or_732_tmp);
  assign and_87_nl = (~ unequal_tmp_4) & equal_tmp_26 & (~ or_732_tmp);
  assign and_89_nl = (~ unequal_tmp_5) & equal_tmp_28 & (~ or_732_tmp);
  assign and_91_nl = (~ unequal_tmp_6) & equal_tmp_30 & (~ or_732_tmp);
  assign and_93_nl = (~ unequal_tmp_7) & equal_tmp_32 & (~ or_732_tmp);
  assign and_95_nl = (~ unequal_tmp_8) & equal_tmp_34 & (~ or_732_tmp);
  assign and_97_nl = (~ unequal_tmp_9) & equal_tmp_36 & (~ or_732_tmp);
  assign and_99_nl = (~ unequal_tmp_10) & equal_tmp_38 & (~ or_732_tmp);
  assign and_101_nl = (~ unequal_tmp_11) & equal_tmp_40 & (~ or_732_tmp);
  assign and_103_nl = (~ unequal_tmp_12) & equal_tmp_42 & (~ or_732_tmp);
  assign and_105_nl = (~ unequal_tmp_13) & equal_tmp_44 & (~ or_732_tmp);
  assign and_107_nl = (~ unequal_tmp_14) & equal_tmp_46 & (~ or_732_tmp);
  assign and_109_nl = (~ unequal_tmp_15) & equal_tmp_48 & (~ or_732_tmp);
  assign and_111_nl = (~ unequal_tmp_16) & equal_tmp_50 & (~ or_732_tmp);
  assign and_203_nl = equal_tmp_52 & (~ or_732_tmp);
  assign mux1h_78_tmp = MUX1HOT_v_5_20_2(({3'b0 , (for_mux_3_nl)}), 5'b11, 5'b100,
      5'b101, 5'b110, 5'b111, 5'b1000, 5'b1001, 5'b1010, 5'b1011, 5'b1100, 5'b1101,
      5'b1110, 5'b1111, 5'b10000, 5'b10001, 5'b10010, 5'b10011, (signext_5_1(nand_17_nl)),
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24, {(and_202_nl) , (and_79_nl) ,
      (and_81_nl) , (and_83_nl) , (and_85_nl) , (and_87_nl) , (and_89_nl) , (and_91_nl)
      , (and_93_nl) , (and_95_nl) , (and_97_nl) , (and_99_nl) , (and_101_nl) , (and_103_nl)
      , (and_105_nl) , (and_107_nl) , (and_109_nl) , (and_111_nl) , (and_203_nl)
      , or_732_tmp});
  assign WRITE_x_idx_6_0_lpi_1_dfm = MUX_v_7_2_2(7'b0000000, WRITE_x_idx_6_0_lpi_2,
      for_unequal_tmp);
  assign unequal_tmp = ~((io_write_dout_0_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_1 = ~((io_write_dout_1_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_2 = ~((io_write_dout_2_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_3 = ~((io_write_dout_3_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_4 = ~((io_write_dout_4_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_5 = ~((io_write_dout_5_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_6 = ~((io_write_dout_6_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_7 = ~((io_write_dout_7_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_8 = ~((io_write_dout_8_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_9 = ~((io_write_dout_9_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_10 = ~((io_write_dout_10_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_11 = ~((io_write_dout_11_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_12 = ~((io_write_dout_12_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_13 = ~((io_write_dout_13_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_14 = ~((io_write_dout_14_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_15 = ~((io_write_dout_15_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign unequal_tmp_16 = ~((io_write_dout_16_copy_ndx_6_0_lpi_1_mx0==7'b1000001));
  assign or_2_tmp_1 = equal_tmp_18 | equal_tmp_20 | equal_tmp_22 | equal_tmp_24 |
      equal_tmp_26 | equal_tmp_28 | equal_tmp_30 | equal_tmp_32 | equal_tmp_34 |
      equal_tmp_36 | equal_tmp_38 | equal_tmp_40 | equal_tmp_42 | equal_tmp_44 |
      equal_tmp_46 | equal_tmp_48 | equal_tmp_50 | equal_tmp_52 | nor_tmp_1;
  assign equal_tmp = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b00010);
  assign equal_tmp_1 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b00011);
  assign equal_tmp_2 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b00100);
  assign equal_tmp_3 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b00101);
  assign equal_tmp_4 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b00110);
  assign equal_tmp_5 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b00111);
  assign equal_tmp_6 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b01000);
  assign equal_tmp_7 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b01001);
  assign equal_tmp_8 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b01010);
  assign equal_tmp_9 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b01011);
  assign equal_tmp_10 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b01100);
  assign equal_tmp_11 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b01101);
  assign equal_tmp_12 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b01110);
  assign equal_tmp_13 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b01111);
  assign equal_tmp_14 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b10000);
  assign equal_tmp_15 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b10001);
  assign equal_tmp_16 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b10010);
  assign nor_tmp = ~(((lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b00001)) | (~((lfst_exit_io_write_dout_17_copy_lpi_1_dfm!=5'b00000)))
      | equal_tmp | equal_tmp_1 | equal_tmp_2 | equal_tmp_3 | equal_tmp_4 | equal_tmp_5
      | equal_tmp_6 | equal_tmp_7 | equal_tmp_8 | equal_tmp_9 | equal_tmp_10 | equal_tmp_11
      | equal_tmp_12 | equal_tmp_13 | equal_tmp_14 | equal_tmp_15 | equal_tmp_16
      | equal_tmp_17);
  assign equal_tmp_17 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm==5'b10011);
  assign nl_WRITE_acc_nl = conv_u2s_6_7(WRITE_x_idx_6_0_sva_1[6:1]) + 7'b1011111;
  assign WRITE_acc_nl = nl_WRITE_acc_nl[6:0];
  assign WRITE_acc_itm_6 = readslicef_7_1_6((WRITE_acc_nl));
  assign nl_WRITE_x_idx_6_0_sva_1 = WRITE_x_idx_6_0_lpi_1_dfm + 7'b1;
  assign WRITE_x_idx_6_0_sva_1 = nl_WRITE_x_idx_6_0_sva_1[6:0];
  assign and_76_rgt = WRITE_for_acc_itm_4_1 & (~ or_1_tmp);
  assign or_1_tmp = equal_tmp | equal_tmp_1 | equal_tmp_2 | equal_tmp_3 | equal_tmp_4
      | equal_tmp_5 | equal_tmp_6 | equal_tmp_7 | equal_tmp_8 | equal_tmp_9 | equal_tmp_10
      | equal_tmp_11 | equal_tmp_12 | equal_tmp_13 | equal_tmp_14 | equal_tmp_15
      | equal_tmp_16 | equal_tmp_17 | nor_tmp;
  assign and_dcpl_19 = ~((mux1h_78_tmp[2:1]!=2'b00));
  assign and_dcpl_20 = ~((mux1h_78_tmp[4:3]!=2'b00));
  assign or_dcpl_8 = (~ main_stage_0_3) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[0]);
  assign or_dcpl_10 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[3]) | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[1]));
  assign or_dcpl_11 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[2]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[4]);
  assign or_dcpl_12 = or_dcpl_11 | or_dcpl_10;
  assign or_dcpl_15 = ~((lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[1]) & main_stage_0_3);
  assign or_dcpl_16 = or_dcpl_15 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[0]);
  assign or_dcpl_17 = or_dcpl_11 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[3]);
  assign or_dcpl_24 = ~(main_stage_0_3 & (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[0]));
  assign or_dcpl_28 = or_dcpl_15 | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[0]));
  assign or_dcpl_36 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[3]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[1]);
  assign or_dcpl_37 = (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[2])) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[4]);
  assign or_dcpl_38 = or_dcpl_37 | or_dcpl_36;
  assign or_dcpl_41 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[1]) | (~ main_stage_0_3);
  assign or_dcpl_42 = or_dcpl_41 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[0]);
  assign or_dcpl_43 = or_dcpl_37 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[3]);
  assign or_dcpl_53 = or_dcpl_41 | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[0]));
  assign or_dcpl_61 = or_dcpl_37 | or_dcpl_10;
  assign or_dcpl_80 = (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[3])) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[1]);
  assign or_dcpl_81 = or_dcpl_11 | or_dcpl_80;
  assign or_dcpl_84 = or_dcpl_11 | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[3]));
  assign or_dcpl_101 = ~((lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[3]) & (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[1]));
  assign or_dcpl_102 = or_dcpl_11 | or_dcpl_101;
  assign or_dcpl_121 = or_dcpl_37 | or_dcpl_80;
  assign or_dcpl_124 = or_dcpl_37 | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[3]));
  assign or_dcpl_141 = or_dcpl_37 | or_dcpl_101;
  assign or_dcpl_160 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[2]) | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[4]));
  assign or_dcpl_161 = or_dcpl_160 | or_dcpl_36;
  assign or_dcpl_164 = or_dcpl_160 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3[3]);
  assign or_dcpl_181 = or_dcpl_160 | or_dcpl_10;
  assign or_dcpl_194 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]);
  assign or_dcpl_195 = or_dcpl_194 | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]));
  assign or_dcpl_196 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]) | (~ main_stage_0_2);
  assign or_dcpl_197 = or_dcpl_196 | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]));
  assign or_dcpl_198 = or_dcpl_197 | or_dcpl_195;
  assign or_dcpl_200 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]) | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]));
  assign or_dcpl_201 = or_dcpl_200 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign or_dcpl_202 = or_dcpl_197 | or_dcpl_201;
  assign or_dcpl_204 = or_dcpl_194 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign or_dcpl_205 = or_dcpl_197 | or_dcpl_204;
  assign or_dcpl_207 = ~((lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]) & (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]));
  assign or_dcpl_208 = or_dcpl_207 | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]));
  assign or_dcpl_210 = (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3])) | (~
      main_stage_0_2) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]);
  assign or_dcpl_211 = or_dcpl_210 | or_dcpl_208;
  assign or_dcpl_213 = (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2])) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]);
  assign or_dcpl_214 = or_dcpl_213 | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]));
  assign or_dcpl_215 = or_dcpl_210 | or_dcpl_214;
  assign or_dcpl_217 = or_dcpl_207 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign or_dcpl_218 = or_dcpl_210 | or_dcpl_217;
  assign or_dcpl_220 = or_dcpl_213 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign or_dcpl_221 = or_dcpl_210 | or_dcpl_220;
  assign or_dcpl_223 = or_dcpl_200 | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]));
  assign or_dcpl_224 = or_dcpl_210 | or_dcpl_223;
  assign or_dcpl_226 = or_dcpl_210 | or_dcpl_195;
  assign or_dcpl_228 = or_dcpl_210 | or_dcpl_201;
  assign or_dcpl_230 = or_dcpl_210 | or_dcpl_204;
  assign or_dcpl_232 = or_dcpl_196 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]);
  assign or_dcpl_233 = or_dcpl_232 | or_dcpl_208;
  assign or_dcpl_235 = or_dcpl_232 | or_dcpl_214;
  assign or_dcpl_237 = or_dcpl_232 | or_dcpl_217;
  assign or_dcpl_239 = or_dcpl_232 | or_dcpl_220;
  assign or_dcpl_241 = or_dcpl_232 | or_dcpl_223;
  assign or_dcpl_243 = or_dcpl_232 | or_dcpl_195;
  assign or_dcpl_246 = or_dcpl_196 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4])
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign or_dcpl_248 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]);
  assign or_dcpl_249 = (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign or_dcpl_250 = or_dcpl_249 | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]);
  assign or_dcpl_251 = or_dcpl_250 | or_dcpl_248;
  assign or_dcpl_253 = or_dcpl_232 | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4:3]!=2'b00);
  assign or_dcpl_256 = or_dcpl_249 | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]));
  assign or_dcpl_257 = or_dcpl_256 | or_dcpl_248;
  assign or_dcpl_260 = or_dcpl_196 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4])
      | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign or_tmp_75 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]) | (~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1]))
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]) | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4])));
  assign or_dcpl_262 = (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign or_dcpl_263 = or_dcpl_262 | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]);
  assign or_dcpl_264 = or_dcpl_263 | or_dcpl_248;
  assign nor_tmp_21 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]) & (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign or_dcpl_267 = or_dcpl_262 | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[0]));
  assign or_dcpl_268 = or_dcpl_267 | or_dcpl_248;
  assign or_dcpl_271 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[2]));
  assign or_dcpl_272 = or_dcpl_250 | or_dcpl_271;
  assign or_dcpl_275 = or_dcpl_256 | or_dcpl_271;
  assign or_dcpl_277 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2:1]!=2'b00);
  assign or_dcpl_278 = (~ main_stage_0_2) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]);
  assign or_dcpl_279 = or_dcpl_278 | or_dcpl_277;
  assign or_tmp_82 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]) | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]));
  assign or_dcpl_281 = or_dcpl_263 | or_dcpl_271;
  assign nor_tmp_23 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]) & (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]);
  assign or_dcpl_284 = or_dcpl_267 | or_dcpl_271;
  assign or_dcpl_286 = or_dcpl_278 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign or_dcpl_289 = or_dcpl_232 | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4:3]!=2'b01);
  assign or_dcpl_293 = or_dcpl_278 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[1]);
  assign nor_tmp_25 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3:2]==2'b11);
  assign or_tmp_90 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]) | (~ nor_tmp_25);
  assign nor_117_nl = ~((~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[1])) | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[3]))
      | (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]) | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]));
  assign mux_tmp_42 = MUX_s_1_2_2((nor_117_nl), (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]),
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign nor_tmp_26 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]) & (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2])
      & (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[3]);
  assign or_dcpl_302 = or_dcpl_196 | or_dcpl_277;
  assign or_tmp_101 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]) | (~ (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]));
  assign nor_tmp_28 = (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[0]) & (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4]);
  assign or_dcpl_307 = or_dcpl_196 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[2]);
  assign or_dcpl_312 = or_dcpl_196 | (lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24[4])
      | (~ (WRITE_for_y_idx_4_0_lpi_1_dfm_st_2[4]));
  assign and_dcpl_28 = ((mux1h_78_tmp[4:1]!=4'b0000)) & main_stage_0_2;
  assign dout_0_rsci_addra_d_pff = io_write_dout_0_copy_ndx_6_0_lpi_1;
  assign dout_0_rsci_dinb_d = dout_0_rsci_dinb_d_reg;
  assign dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_1_rsci_addra_d_pff = io_write_dout_1_copy_ndx_6_0_lpi_1;
  assign dout_1_rsci_dinb_d = dout_1_rsci_dinb_d_reg;
  assign dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_2_rsci_addra_d_pff = io_write_dout_2_copy_ndx_6_0_lpi_1;
  assign dout_2_rsci_dinb_d = dout_2_rsci_dinb_d_reg;
  assign dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_3_rsci_addra_d_pff = io_write_dout_3_copy_ndx_6_0_lpi_1;
  assign dout_3_rsci_dinb_d = dout_3_rsci_dinb_d_reg;
  assign dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_4_rsci_addra_d_pff = io_write_dout_4_copy_ndx_6_0_lpi_1;
  assign dout_4_rsci_dinb_d = dout_4_rsci_dinb_d_reg;
  assign dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_5_rsci_addra_d_pff = io_write_dout_5_copy_ndx_6_0_lpi_1;
  assign dout_5_rsci_dinb_d = dout_5_rsci_dinb_d_reg;
  assign dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_6_rsci_addra_d_pff = io_write_dout_6_copy_ndx_6_0_lpi_1;
  assign dout_6_rsci_dinb_d = dout_6_rsci_dinb_d_reg;
  assign dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_7_rsci_addra_d_pff = io_write_dout_7_copy_ndx_6_0_lpi_1;
  assign dout_7_rsci_dinb_d = dout_7_rsci_dinb_d_reg;
  assign dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_8_rsci_addra_d_pff = io_write_dout_8_copy_ndx_6_0_lpi_1;
  assign dout_8_rsci_dinb_d = dout_8_rsci_dinb_d_reg;
  assign dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_9_rsci_addra_d_pff = io_write_dout_9_copy_ndx_6_0_lpi_1;
  assign dout_9_rsci_dinb_d = dout_9_rsci_dinb_d_reg;
  assign dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_10_rsci_addra_d_pff = io_write_dout_10_copy_ndx_6_0_lpi_1;
  assign dout_10_rsci_dinb_d = dout_10_rsci_dinb_d_reg;
  assign dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_11_rsci_addra_d_pff = io_write_dout_11_copy_ndx_6_0_lpi_1;
  assign dout_11_rsci_dinb_d = dout_11_rsci_dinb_d_reg;
  assign dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_12_rsci_addra_d_pff = io_write_dout_12_copy_ndx_6_0_lpi_1;
  assign dout_12_rsci_dinb_d = dout_12_rsci_dinb_d_reg;
  assign dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_13_rsci_addra_d_pff = io_write_dout_13_copy_ndx_6_0_lpi_1;
  assign dout_13_rsci_dinb_d = dout_13_rsci_dinb_d_reg;
  assign dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_14_rsci_addra_d_pff = io_write_dout_14_copy_ndx_6_0_lpi_1;
  assign dout_14_rsci_dinb_d = dout_14_rsci_dinb_d_reg;
  assign dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_15_rsci_addra_d_pff = io_write_dout_15_copy_ndx_6_0_lpi_1;
  assign dout_15_rsci_dinb_d = dout_15_rsci_dinb_d_reg;
  assign dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_16_rsci_addra_d_pff = io_write_dout_16_copy_ndx_6_0_lpi_1;
  assign dout_16_rsci_dinb_d = dout_16_rsci_dinb_d_reg;
  assign dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_17_rsci_addra_d_pff = io_write_dout_17_copy_ndx_6_0_lpi_1;
  assign dout_17_rsci_dinb_d = dout_17_rsci_dinb_d_reg;
  assign dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_0_data_rsci_addra_d = tmp_0_data_rsci_addra_d_reg;
  assign tmp_0_data_rsci_addrb_d = tmp_0_data_rsci_addrb_d_reg;
  assign tmp_0_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_1_data_rsci_addra_d = tmp_1_data_rsci_addra_d_reg;
  assign tmp_1_data_rsci_addrb_d = tmp_1_data_rsci_addrb_d_reg;
  assign tmp_1_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_2_data_rsci_addra_d = tmp_2_data_rsci_addra_d_reg;
  assign tmp_2_data_rsci_addrb_d = tmp_2_data_rsci_addrb_d_reg;
  assign tmp_2_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_3_data_rsci_addra_d = tmp_3_data_rsci_addra_d_reg;
  assign tmp_3_data_rsci_addrb_d = tmp_3_data_rsci_addrb_d_reg;
  assign tmp_3_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_4_data_rsci_addra_d = tmp_4_data_rsci_addra_d_reg;
  assign tmp_4_data_rsci_addrb_d = tmp_4_data_rsci_addrb_d_reg;
  assign tmp_4_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_5_data_rsci_addra_d = tmp_5_data_rsci_addra_d_reg;
  assign tmp_5_data_rsci_addrb_d = tmp_5_data_rsci_addrb_d_reg;
  assign tmp_5_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_6_data_rsci_addra_d = tmp_6_data_rsci_addra_d_reg;
  assign tmp_6_data_rsci_addrb_d = tmp_6_data_rsci_addrb_d_reg;
  assign tmp_6_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_7_data_rsci_addra_d = tmp_7_data_rsci_addra_d_reg;
  assign tmp_7_data_rsci_addrb_d = tmp_7_data_rsci_addrb_d_reg;
  assign tmp_7_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_8_data_rsci_addra_d = tmp_8_data_rsci_addra_d_reg;
  assign tmp_8_data_rsci_addrb_d = tmp_8_data_rsci_addrb_d_reg;
  assign tmp_8_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_9_data_rsci_addra_d = tmp_9_data_rsci_addra_d_reg;
  assign tmp_9_data_rsci_addrb_d = tmp_9_data_rsci_addrb_d_reg;
  assign tmp_9_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_10_data_rsci_addra_d = tmp_10_data_rsci_addra_d_reg;
  assign tmp_10_data_rsci_addrb_d = tmp_10_data_rsci_addrb_d_reg;
  assign tmp_10_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_11_data_rsci_addra_d = tmp_11_data_rsci_addra_d_reg;
  assign tmp_11_data_rsci_addrb_d = tmp_11_data_rsci_addrb_d_reg;
  assign tmp_11_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_12_data_rsci_addra_d = tmp_12_data_rsci_addra_d_reg;
  assign tmp_12_data_rsci_addrb_d = tmp_12_data_rsci_addrb_d_reg;
  assign tmp_12_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_13_data_rsci_addra_d = tmp_13_data_rsci_addra_d_reg;
  assign tmp_13_data_rsci_addrb_d = tmp_13_data_rsci_addrb_d_reg;
  assign tmp_13_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_14_data_rsci_addra_d = tmp_14_data_rsci_addra_d_reg;
  assign tmp_14_data_rsci_addrb_d = tmp_14_data_rsci_addrb_d_reg;
  assign tmp_14_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_15_data_rsci_addra_d = tmp_15_data_rsci_addra_d_reg;
  assign tmp_15_data_rsci_addrb_d = tmp_15_data_rsci_addrb_d_reg;
  assign tmp_15_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_16_data_rsci_addra_d = tmp_16_data_rsci_addra_d_reg;
  assign tmp_16_data_rsci_addrb_d = tmp_16_data_rsci_addrb_d_reg;
  assign tmp_16_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign tmp_17_data_rsci_addra_d = tmp_17_data_rsci_addra_d_reg;
  assign tmp_17_data_rsci_addrb_d = tmp_17_data_rsci_addrb_d_reg;
  assign tmp_17_data_rsci_dinb_d = {{48{din_rsci_d_mxwt[15]}}, din_rsci_d_mxwt};
  assign tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      reg_dout_0_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_1_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_2_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_3_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_4_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_5_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_6_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_7_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_8_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_9_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_10_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_11_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_12_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_13_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_14_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_15_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_16_rsc_rls_obj_iswt0_cse <= 1'b0;
      reg_dout_17_rsc_rls_obj_iswt0_cse <= 1'b0;
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24 <= 5'b0;
      reg_dout_17_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_16_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_15_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_14_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_13_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_12_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_11_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_10_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_9_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_8_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_7_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_6_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_5_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_4_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_3_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_2_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_1_rsc_req_obj_oswt_cse <= 1'b0;
      nor_dfs_3 <= 1'b0;
      equal_tmp_72 <= 1'b0;
      equal_tmp_73 <= 1'b0;
      equal_tmp_74 <= 1'b0;
      equal_tmp_75 <= 1'b0;
      equal_tmp_76 <= 1'b0;
      equal_tmp_77 <= 1'b0;
      equal_tmp_78 <= 1'b0;
      equal_tmp_79 <= 1'b0;
      equal_tmp_80 <= 1'b0;
      equal_tmp_81 <= 1'b0;
      equal_tmp_82 <= 1'b0;
      equal_tmp_83 <= 1'b0;
      equal_tmp_84 <= 1'b0;
      equal_tmp_85 <= 1'b0;
      equal_tmp_86 <= 1'b0;
      equal_tmp_87 <= 1'b0;
      nor_tmp_30 <= 1'b0;
      equal_tmp_88 <= 1'b0;
      equal_tmp_89 <= 1'b0;
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3 <= 5'b0;
      reg_tmp_0_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_1_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_2_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_3_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_4_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_5_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_6_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_7_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_8_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_9_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_10_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_11_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_12_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_13_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_14_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_15_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_16_data_rsci_oswt_cse <= 1'b0;
      reg_tmp_17_data_rsci_oswt_cse <= 1'b0;
      reg_dout_0_rsc_req_obj_oswt_cse <= 1'b0;
      reg_din_rsci_oswt_cse <= 1'b0;
      lfst_exit_WRITE_lpi_1 <= 1'b0;
      WRITE_x_idx_6_0_lpi_1_dfm_5 <= 7'b0;
      WRITE_for_y_idx_4_0_lpi_1_dfm_st_2 <= 5'b0;
      exit_WRITE_lpi_1_dfm_4 <= 1'b0;
      WRITE_for_slc_WRITE_for_acc_4_svs_2 <= 1'b0;
      equal_tmp_18 <= 1'b0;
      equal_tmp_20 <= 1'b0;
      equal_tmp_22 <= 1'b0;
      equal_tmp_24 <= 1'b0;
      equal_tmp_26 <= 1'b0;
      equal_tmp_28 <= 1'b0;
      equal_tmp_30 <= 1'b0;
      equal_tmp_32 <= 1'b0;
      equal_tmp_34 <= 1'b0;
      equal_tmp_36 <= 1'b0;
      equal_tmp_38 <= 1'b0;
      equal_tmp_40 <= 1'b0;
      equal_tmp_42 <= 1'b0;
      equal_tmp_44 <= 1'b0;
      equal_tmp_46 <= 1'b0;
      equal_tmp_48 <= 1'b0;
      equal_tmp_50 <= 1'b0;
      nor_tmp_1 <= 1'b0;
      equal_tmp_52 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_dout_0_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_12 | or_dcpl_8 | (io_write_dout_0_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_1_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_12 | or_dcpl_24 | (io_write_dout_1_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_2_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_38 | or_dcpl_8 | (io_write_dout_2_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_3_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_38 | or_dcpl_24 | (io_write_dout_3_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_4_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_61 | or_dcpl_8 | (io_write_dout_4_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_5_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_61 | or_dcpl_24 | (io_write_dout_5_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_6_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_81 | or_dcpl_8 | (io_write_dout_6_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_7_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_81 | or_dcpl_24 | (io_write_dout_7_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_8_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_102 | or_dcpl_8 | (io_write_dout_8_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_9_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_102 | or_dcpl_24 | (io_write_dout_9_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_10_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_121 | or_dcpl_8 | (io_write_dout_10_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_11_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_121 | or_dcpl_24 | (io_write_dout_11_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_12_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_141 | or_dcpl_8 | (io_write_dout_12_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_13_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_141 | or_dcpl_24 | (io_write_dout_13_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_14_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_161 | or_dcpl_8 | (io_write_dout_14_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_15_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_161 | or_dcpl_24 | (io_write_dout_15_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_16_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_181 | or_dcpl_8 | (io_write_dout_16_copy_ndx_6_0_lpi_1!=7'b1000001));
      reg_dout_17_rsc_rls_obj_iswt0_cse <= ~(or_dcpl_181 | or_dcpl_24 | (io_write_dout_17_copy_ndx_6_0_lpi_1!=7'b1000001));
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24 <= lfst_exit_io_write_dout_17_copy_lpi_1_dfm;
      reg_dout_17_rsc_req_obj_oswt_cse <= ~((mux_132_nl) | or_dcpl_198);
      reg_dout_16_rsc_req_obj_oswt_cse <= ~((mux_133_nl) | or_dcpl_202);
      reg_dout_15_rsc_req_obj_oswt_cse <= ~((mux_134_nl) | or_dcpl_205);
      reg_dout_14_rsc_req_obj_oswt_cse <= ~((mux_135_nl) | or_dcpl_211);
      reg_dout_13_rsc_req_obj_oswt_cse <= ~((mux_136_nl) | or_dcpl_215);
      reg_dout_12_rsc_req_obj_oswt_cse <= ~((mux_137_nl) | or_dcpl_218);
      reg_dout_11_rsc_req_obj_oswt_cse <= ~((mux_138_nl) | or_dcpl_221);
      reg_dout_10_rsc_req_obj_oswt_cse <= ~((mux_139_nl) | or_dcpl_224);
      reg_dout_9_rsc_req_obj_oswt_cse <= ~((mux_140_nl) | or_dcpl_226);
      reg_dout_8_rsc_req_obj_oswt_cse <= ~((mux_141_nl) | or_dcpl_228);
      reg_dout_7_rsc_req_obj_oswt_cse <= ~((mux_142_nl) | or_dcpl_230);
      reg_dout_6_rsc_req_obj_oswt_cse <= ~((mux_143_nl) | or_dcpl_233);
      reg_dout_5_rsc_req_obj_oswt_cse <= ~((mux_144_nl) | or_dcpl_235);
      reg_dout_4_rsc_req_obj_oswt_cse <= ~((mux_145_nl) | or_dcpl_237);
      reg_dout_3_rsc_req_obj_oswt_cse <= ~((mux_146_nl) | or_dcpl_239);
      reg_dout_2_rsc_req_obj_oswt_cse <= ~((mux_147_nl) | or_dcpl_241);
      reg_dout_1_rsc_req_obj_oswt_cse <= ~((mux_148_nl) | or_dcpl_243);
      nor_dfs_3 <= nor_19_tmp;
      equal_tmp_72 <= equal_tmp_18;
      equal_tmp_73 <= equal_tmp_20;
      equal_tmp_74 <= equal_tmp_22;
      equal_tmp_75 <= equal_tmp_24;
      equal_tmp_76 <= equal_tmp_26;
      equal_tmp_77 <= equal_tmp_28;
      equal_tmp_78 <= equal_tmp_30;
      equal_tmp_79 <= equal_tmp_32;
      equal_tmp_80 <= equal_tmp_34;
      equal_tmp_81 <= equal_tmp_36;
      equal_tmp_82 <= equal_tmp_38;
      equal_tmp_83 <= equal_tmp_40;
      equal_tmp_84 <= equal_tmp_42;
      equal_tmp_85 <= equal_tmp_44;
      equal_tmp_86 <= equal_tmp_46;
      equal_tmp_87 <= equal_tmp_48;
      nor_tmp_30 <= nor_tmp_1;
      equal_tmp_88 <= equal_tmp_50;
      equal_tmp_89 <= equal_tmp_52;
      lfst_exit_io_write_dout_17_copy_lpi_1_dfm_st_3 <= lfst_exit_io_write_dout_17_copy_lpi_1_dfm_24;
      reg_tmp_0_data_rsci_oswt_cse <= WRITE_for_if_nor_rmff;
      reg_tmp_1_data_rsci_oswt_cse <= WRITE_for_else_if_nor_rmff;
      reg_tmp_2_data_rsci_oswt_cse <= WRITE_for_else_else_if_nor_rmff;
      reg_tmp_3_data_rsci_oswt_cse <= WRITE_for_else_else_else_if_nor_rmff;
      reg_tmp_4_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_if_nor_rmff;
      reg_tmp_5_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_if_nor_rmff;
      reg_tmp_6_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_7_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_8_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_9_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_10_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_11_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_12_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_13_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_14_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_15_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_16_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
      reg_tmp_17_data_rsci_oswt_cse <= WRITE_for_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_else_if_nor_rmff;
      reg_dout_0_rsc_req_obj_oswt_cse <= ~(or_dcpl_232 | or_dcpl_277 | (~ exit_WRITE_lpi_1_dfm_4));
      reg_din_rsci_oswt_cse <= ~ and_dcpl_28;
      lfst_exit_WRITE_lpi_1 <= lfst_exit_WRITE_lpi_1_mx0;
      WRITE_x_idx_6_0_lpi_1_dfm_5 <= WRITE_x_idx_6_0_lpi_1_dfm;
      WRITE_for_y_idx_4_0_lpi_1_dfm_st_2 <= WRITE_for_y_idx_4_0_lpi_1_dfm;
      exit_WRITE_lpi_1_dfm_4 <= ~(WRITE_acc_itm_6 | WRITE_for_acc_itm_4_1);
      WRITE_for_slc_WRITE_for_acc_4_svs_2 <= WRITE_for_acc_itm_4_1;
      equal_tmp_18 <= equal_tmp;
      equal_tmp_20 <= equal_tmp_1;
      equal_tmp_22 <= equal_tmp_2;
      equal_tmp_24 <= equal_tmp_3;
      equal_tmp_26 <= equal_tmp_4;
      equal_tmp_28 <= equal_tmp_5;
      equal_tmp_30 <= equal_tmp_6;
      equal_tmp_32 <= equal_tmp_7;
      equal_tmp_34 <= equal_tmp_8;
      equal_tmp_36 <= equal_tmp_9;
      equal_tmp_38 <= equal_tmp_10;
      equal_tmp_40 <= equal_tmp_11;
      equal_tmp_42 <= equal_tmp_12;
      equal_tmp_44 <= equal_tmp_13;
      equal_tmp_46 <= equal_tmp_14;
      equal_tmp_48 <= equal_tmp_15;
      equal_tmp_50 <= equal_tmp_16;
      nor_tmp_1 <= nor_tmp;
      equal_tmp_52 <= equal_tmp_17;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_0_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (or_3_tmp | equal_tmp_72 | nor_dfs_3 | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_0_copy_ndx_6_0_lpi_1 <= io_write_dout_0_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_1_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_73 | equal_tmp_72 | or_4_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_1_copy_ndx_6_0_lpi_1 <= io_write_dout_1_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_2_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_74 | equal_tmp_73 | or_5_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_2_copy_ndx_6_0_lpi_1 <= io_write_dout_2_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_3_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_75 | equal_tmp_74 | or_6_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_3_copy_ndx_6_0_lpi_1 <= io_write_dout_3_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_4_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_76 | equal_tmp_75 | or_7_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_4_copy_ndx_6_0_lpi_1 <= io_write_dout_4_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_5_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_77 | equal_tmp_76 | or_8_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_5_copy_ndx_6_0_lpi_1 <= io_write_dout_5_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_6_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_78 | equal_tmp_77 | or_9_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_6_copy_ndx_6_0_lpi_1 <= io_write_dout_6_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_7_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_79 | equal_tmp_78 | or_10_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_7_copy_ndx_6_0_lpi_1 <= io_write_dout_7_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_8_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_80 | equal_tmp_79 | or_11_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_8_copy_ndx_6_0_lpi_1 <= io_write_dout_8_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_9_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_81 | equal_tmp_80 | or_12_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_9_copy_ndx_6_0_lpi_1 <= io_write_dout_9_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_10_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_82 | equal_tmp_81 | or_13_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_10_copy_ndx_6_0_lpi_1 <= io_write_dout_10_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_11_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_83 | equal_tmp_82 | or_14_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_11_copy_ndx_6_0_lpi_1 <= io_write_dout_11_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_12_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_84 | equal_tmp_83 | or_15_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_12_copy_ndx_6_0_lpi_1 <= io_write_dout_12_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_13_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_85 | equal_tmp_84 | or_16_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_13_copy_ndx_6_0_lpi_1 <= io_write_dout_13_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_14_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_86 | equal_tmp_85 | or_17_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_14_copy_ndx_6_0_lpi_1 <= io_write_dout_14_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_15_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_87 | equal_tmp_86 | or_18_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_15_copy_ndx_6_0_lpi_1 <= io_write_dout_15_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_16_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_88 | equal_tmp_87 | or_19_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_16_copy_ndx_6_0_lpi_1 <= io_write_dout_16_copy_ndx_6_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_17_copy_ndx_6_0_lpi_1 <= 7'b0;
    end
    else if ( (equal_tmp_89 | equal_tmp_88 | or_20_tmp | (~ main_stage_0_3)) & core_wen
        ) begin
      io_write_dout_17_copy_ndx_6_0_lpi_1 <= mux_53_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_17_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_16_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_206_cse ) begin
      io_write_dout_17_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, mux_53_tmp,
          unequal_tmp_16);
      io_write_dout_16_copy_ndx_6_0_sva_4 <= nl_io_write_dout_16_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_17_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( core_wen & main_stage_0_2 & equal_tmp_52 ) begin
      io_write_dout_17_copy_ndx_6_0_sva_4 <= nl_io_write_dout_17_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_16_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_15_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_208_cse ) begin
      io_write_dout_16_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_16_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_15);
      io_write_dout_15_copy_ndx_6_0_sva_4 <= nl_io_write_dout_15_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_15_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_14_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_210_cse ) begin
      io_write_dout_15_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_15_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_14);
      io_write_dout_14_copy_ndx_6_0_sva_4 <= nl_io_write_dout_14_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_14_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_13_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_212_cse ) begin
      io_write_dout_14_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_14_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_13);
      io_write_dout_13_copy_ndx_6_0_sva_4 <= nl_io_write_dout_13_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_13_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_12_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_214_cse ) begin
      io_write_dout_13_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_13_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_12);
      io_write_dout_12_copy_ndx_6_0_sva_4 <= nl_io_write_dout_12_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_12_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_11_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_216_cse ) begin
      io_write_dout_12_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_12_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_11);
      io_write_dout_11_copy_ndx_6_0_sva_4 <= nl_io_write_dout_11_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_11_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_10_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_218_cse ) begin
      io_write_dout_11_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_11_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_10);
      io_write_dout_10_copy_ndx_6_0_sva_4 <= nl_io_write_dout_10_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_10_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_9_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_220_cse ) begin
      io_write_dout_10_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_10_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_9);
      io_write_dout_9_copy_ndx_6_0_sva_4 <= nl_io_write_dout_9_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_9_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_8_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_222_cse ) begin
      io_write_dout_9_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_9_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_8);
      io_write_dout_8_copy_ndx_6_0_sva_4 <= nl_io_write_dout_8_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_8_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_7_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_224_cse ) begin
      io_write_dout_8_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_8_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_7);
      io_write_dout_7_copy_ndx_6_0_sva_4 <= nl_io_write_dout_7_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_7_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_6_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_226_cse ) begin
      io_write_dout_7_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_7_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_6);
      io_write_dout_6_copy_ndx_6_0_sva_4 <= nl_io_write_dout_6_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_6_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_5_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_228_cse ) begin
      io_write_dout_6_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_6_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_5);
      io_write_dout_5_copy_ndx_6_0_sva_4 <= nl_io_write_dout_5_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_5_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_4_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_230_cse ) begin
      io_write_dout_5_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_5_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_4);
      io_write_dout_4_copy_ndx_6_0_sva_4 <= nl_io_write_dout_4_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_4_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_3_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_232_cse ) begin
      io_write_dout_4_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_4_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_3);
      io_write_dout_3_copy_ndx_6_0_sva_4 <= nl_io_write_dout_3_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_3_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_2_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_234_cse ) begin
      io_write_dout_3_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_3_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_2);
      io_write_dout_2_copy_ndx_6_0_sva_4 <= nl_io_write_dout_2_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_2_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_1_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_236_cse ) begin
      io_write_dout_2_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_2_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp_1);
      io_write_dout_1_copy_ndx_6_0_sva_4 <= nl_io_write_dout_1_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_1_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
      io_write_dout_0_copy_ndx_6_0_sva_4 <= 7'b0;
    end
    else if ( and_238_cse ) begin
      io_write_dout_1_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_1_copy_ndx_6_0_lpi_1_mx0,
          unequal_tmp);
      io_write_dout_0_copy_ndx_6_0_sva_4 <= nl_io_write_dout_0_copy_ndx_6_0_sva_4[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      io_write_dout_0_copy_ndx_6_0_lpi_1_dfm_4 <= 7'b0;
    end
    else if ( core_wen & main_stage_0_2 & nor_19_tmp ) begin
      io_write_dout_0_copy_ndx_6_0_lpi_1_dfm_4 <= MUX_v_7_2_2(7'b0000000, io_write_dout_0_copy_ndx_6_0_lpi_1_mx0,
          (WRITE_not_8_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      WRITE_for_y_idx_4_0_lpi_3 <= 5'b0;
    end
    else if ( core_wen & main_stage_0_2 & mux_130_cse ) begin
      WRITE_for_y_idx_4_0_lpi_3 <= mux1h_77_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      WRITE_for_y_idx_slc_WRITE_for_y_idx_4_0_0_itm_3 <= 1'b0;
    end
    else if ( core_wen & mux_130_cse & and_dcpl_20 & and_dcpl_19 & main_stage_0_2
        & (mux1h_78_tmp[0]) & (mux1h_77_tmp[4]) ) begin
      WRITE_for_y_idx_slc_WRITE_for_y_idx_4_0_0_itm_3 <= WRITE_for_y_idx_4_0_lpi_1_dfm[0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      WRITE_for_y_idx_4_0_sva_6 <= 5'b0;
    end
    else if ( core_wen & (~((~(and_dcpl_20 & and_dcpl_19)) & main_stage_0_2)) & WRITE_for_acc_itm_4_1
        ) begin
      WRITE_for_y_idx_4_0_sva_6 <= WRITE_for_y_idx_4_0_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exit_WRITE_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_28 | WRITE_for_acc_itm_4_1)) ) begin
      exit_WRITE_sva_2 <= ~ WRITE_acc_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      WRITE_x_idx_6_0_lpi_2 <= 7'b0;
    end
    else if ( core_wen & ((~(WRITE_for_acc_itm_4_1 | or_1_tmp)) | and_76_rgt) ) begin
      WRITE_x_idx_6_0_lpi_2 <= MUX_v_7_2_2(WRITE_x_idx_6_0_sva_1, WRITE_x_idx_6_0_lpi_1_dfm,
          and_76_rgt);
    end
  end
  assign and_141_nl = main_stage_0_3 & ((mux1h_19_tmp!=7'b1000001));
  assign or_245_nl = (~ main_stage_0_3) | (mux1h_19_tmp!=7'b1000001);
  assign nor_76_nl = ~((io_write_dout_16_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_132_nl = MUX_s_1_2_2((or_245_nl), (and_141_nl), nor_76_nl);
  assign and_142_nl = main_stage_0_3 & ((mux1h_18_tmp!=7'b1000001));
  assign or_253_nl = (~ main_stage_0_3) | (mux1h_18_tmp!=7'b1000001);
  assign nor_77_nl = ~((io_write_dout_15_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_133_nl = MUX_s_1_2_2((or_253_nl), (and_142_nl), nor_77_nl);
  assign and_143_nl = main_stage_0_3 & ((mux1h_17_tmp!=7'b1000001));
  assign or_260_nl = (~ main_stage_0_3) | (mux1h_17_tmp!=7'b1000001);
  assign nor_78_nl = ~((io_write_dout_14_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_134_nl = MUX_s_1_2_2((or_260_nl), (and_143_nl), nor_78_nl);
  assign and_144_nl = main_stage_0_3 & ((mux1h_16_tmp!=7'b1000001));
  assign or_270_nl = (~ main_stage_0_3) | (mux1h_16_tmp!=7'b1000001);
  assign nor_79_nl = ~((io_write_dout_13_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_135_nl = MUX_s_1_2_2((or_270_nl), (and_144_nl), nor_79_nl);
  assign and_145_nl = main_stage_0_3 & ((mux1h_15_tmp!=7'b1000001));
  assign or_278_nl = (~ main_stage_0_3) | (mux1h_15_tmp!=7'b1000001);
  assign nor_80_nl = ~((io_write_dout_12_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_136_nl = MUX_s_1_2_2((or_278_nl), (and_145_nl), nor_80_nl);
  assign and_146_nl = main_stage_0_3 & ((mux1h_14_tmp!=7'b1000001));
  assign or_285_nl = (~ main_stage_0_3) | (mux1h_14_tmp!=7'b1000001);
  assign nor_81_nl = ~((io_write_dout_11_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_137_nl = MUX_s_1_2_2((or_285_nl), (and_146_nl), nor_81_nl);
  assign and_147_nl = main_stage_0_3 & ((mux1h_13_tmp!=7'b1000001));
  assign or_292_nl = (~ main_stage_0_3) | (mux1h_13_tmp!=7'b1000001);
  assign nor_82_nl = ~((io_write_dout_10_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_138_nl = MUX_s_1_2_2((or_292_nl), (and_147_nl), nor_82_nl);
  assign and_148_nl = main_stage_0_3 & ((mux1h_12_tmp!=7'b1000001));
  assign or_299_nl = (~ main_stage_0_3) | (mux1h_12_tmp!=7'b1000001);
  assign nor_83_nl = ~((io_write_dout_9_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_139_nl = MUX_s_1_2_2((or_299_nl), (and_148_nl), nor_83_nl);
  assign and_149_nl = main_stage_0_3 & ((mux1h_11_tmp!=7'b1000001));
  assign or_305_nl = (~ main_stage_0_3) | (mux1h_11_tmp!=7'b1000001);
  assign nor_84_nl = ~((io_write_dout_8_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_140_nl = MUX_s_1_2_2((or_305_nl), (and_149_nl), nor_84_nl);
  assign and_150_nl = main_stage_0_3 & ((mux1h_10_tmp!=7'b1000001));
  assign or_311_nl = (~ main_stage_0_3) | (mux1h_10_tmp!=7'b1000001);
  assign nor_85_nl = ~((io_write_dout_7_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_141_nl = MUX_s_1_2_2((or_311_nl), (and_150_nl), nor_85_nl);
  assign and_151_nl = main_stage_0_3 & ((mux1h_9_tmp!=7'b1000001));
  assign or_317_nl = (~ main_stage_0_3) | (mux1h_9_tmp!=7'b1000001);
  assign nor_86_nl = ~((io_write_dout_6_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_142_nl = MUX_s_1_2_2((or_317_nl), (and_151_nl), nor_86_nl);
  assign and_152_nl = main_stage_0_3 & ((mux1h_8_tmp!=7'b1000001));
  assign or_324_nl = (~ main_stage_0_3) | (mux1h_8_tmp!=7'b1000001);
  assign nor_87_nl = ~((io_write_dout_5_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_143_nl = MUX_s_1_2_2((or_324_nl), (and_152_nl), nor_87_nl);
  assign and_153_nl = main_stage_0_3 & ((mux1h_7_tmp!=7'b1000001));
  assign or_330_nl = (~ main_stage_0_3) | (mux1h_7_tmp!=7'b1000001);
  assign nor_88_nl = ~((io_write_dout_4_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_144_nl = MUX_s_1_2_2((or_330_nl), (and_153_nl), nor_88_nl);
  assign and_154_nl = main_stage_0_3 & ((mux1h_6_tmp!=7'b1000001));
  assign or_336_nl = (~ main_stage_0_3) | (mux1h_6_tmp!=7'b1000001);
  assign nor_89_nl = ~((io_write_dout_3_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_145_nl = MUX_s_1_2_2((or_336_nl), (and_154_nl), nor_89_nl);
  assign and_155_nl = main_stage_0_3 & ((mux1h_5_tmp!=7'b1000001));
  assign or_342_nl = (~ main_stage_0_3) | (mux1h_5_tmp!=7'b1000001);
  assign nor_90_nl = ~((io_write_dout_2_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_146_nl = MUX_s_1_2_2((or_342_nl), (and_155_nl), nor_90_nl);
  assign and_156_nl = main_stage_0_3 & ((mux1h_4_tmp!=7'b1000001));
  assign or_348_nl = (~ main_stage_0_3) | (mux1h_4_tmp!=7'b1000001);
  assign nor_91_nl = ~((io_write_dout_1_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_147_nl = MUX_s_1_2_2((or_348_nl), (and_156_nl), nor_91_nl);
  assign and_157_nl = main_stage_0_3 & ((mux1h_3_tmp!=7'b1000001));
  assign or_354_nl = (~ main_stage_0_3) | (mux1h_3_tmp!=7'b1000001);
  assign nor_92_nl = ~((io_write_dout_0_copy_ndx_6_0_lpi_1!=7'b1000001));
  assign mux_148_nl = MUX_s_1_2_2((or_354_nl), (and_157_nl), nor_92_nl);
  assign nl_io_write_dout_16_copy_ndx_6_0_sva_4  = io_write_dout_16_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_17_copy_ndx_6_0_sva_4  = mux_53_tmp + 7'b1;
  assign nl_io_write_dout_15_copy_ndx_6_0_sva_4  = io_write_dout_15_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_14_copy_ndx_6_0_sva_4  = io_write_dout_14_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_13_copy_ndx_6_0_sva_4  = io_write_dout_13_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_12_copy_ndx_6_0_sva_4  = io_write_dout_12_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_11_copy_ndx_6_0_sva_4  = io_write_dout_11_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_10_copy_ndx_6_0_sva_4  = io_write_dout_10_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_9_copy_ndx_6_0_sva_4  = io_write_dout_9_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_8_copy_ndx_6_0_sva_4  = io_write_dout_8_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_7_copy_ndx_6_0_sva_4  = io_write_dout_7_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_6_copy_ndx_6_0_sva_4  = io_write_dout_6_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_5_copy_ndx_6_0_sva_4  = io_write_dout_5_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_4_copy_ndx_6_0_sva_4  = io_write_dout_4_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_3_copy_ndx_6_0_sva_4  = io_write_dout_3_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_2_copy_ndx_6_0_sva_4  = io_write_dout_2_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_1_copy_ndx_6_0_sva_4  = io_write_dout_1_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign nl_io_write_dout_0_copy_ndx_6_0_sva_4  = io_write_dout_0_copy_ndx_6_0_lpi_1_mx0
      + 7'b1;
  assign WRITE_not_8_nl = ~ exit_WRITE_lpi_1_dfm_4;

  function [4:0] MUX1HOT_v_5_20_2;
    input [4:0] input_19;
    input [4:0] input_18;
    input [4:0] input_17;
    input [4:0] input_16;
    input [4:0] input_15;
    input [4:0] input_14;
    input [4:0] input_13;
    input [4:0] input_12;
    input [4:0] input_11;
    input [4:0] input_10;
    input [4:0] input_9;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [19:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    result = result | ( input_4 & {5{sel[4]}});
    result = result | ( input_5 & {5{sel[5]}});
    result = result | ( input_6 & {5{sel[6]}});
    result = result | ( input_7 & {5{sel[7]}});
    result = result | ( input_8 & {5{sel[8]}});
    result = result | ( input_9 & {5{sel[9]}});
    result = result | ( input_10 & {5{sel[10]}});
    result = result | ( input_11 & {5{sel[11]}});
    result = result | ( input_12 & {5{sel[12]}});
    result = result | ( input_13 & {5{sel[13]}});
    result = result | ( input_14 & {5{sel[14]}});
    result = result | ( input_15 & {5{sel[15]}});
    result = result | ( input_16 & {5{sel[16]}});
    result = result | ( input_17 & {5{sel[17]}});
    result = result | ( input_18 & {5{sel[18]}});
    result = result | ( input_19 & {5{sel[19]}});
    MUX1HOT_v_5_20_2 = result;
  end
  endfunction


  function [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function [4:0] signext_5_1;
    input [0:0] vector;
  begin
    signext_5_1= {{4{vector[0]}}, vector};
  end
  endfunction


  function  [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function  [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core (
  clk, rst, din_0_rsc_req_vz, din_0_rsc_rls_lz, din_1_rsc_req_vz, din_1_rsc_rls_lz,
      din_2_rsc_req_vz, din_2_rsc_rls_lz, din_3_rsc_req_vz, din_3_rsc_rls_lz, din_4_rsc_req_vz,
      din_4_rsc_rls_lz, din_5_rsc_req_vz, din_5_rsc_rls_lz, din_6_rsc_req_vz, din_6_rsc_rls_lz,
      din_7_rsc_req_vz, din_7_rsc_rls_lz, din_8_rsc_req_vz, din_8_rsc_rls_lz, din_9_rsc_req_vz,
      din_9_rsc_rls_lz, din_10_rsc_req_vz, din_10_rsc_rls_lz, din_11_rsc_req_vz,
      din_11_rsc_rls_lz, din_12_rsc_req_vz, din_12_rsc_rls_lz, din_13_rsc_req_vz,
      din_13_rsc_rls_lz, din_14_rsc_req_vz, din_14_rsc_rls_lz, din_15_rsc_req_vz,
      din_15_rsc_rls_lz, din_16_rsc_req_vz, din_16_rsc_rls_lz, din_17_rsc_req_vz,
      din_17_rsc_rls_lz, dout_rsc_z, dout_rsc_vz, dout_rsc_lz, din_0_rsci_douta_d,
      din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_1_rsci_douta_d, din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_2_rsci_douta_d, din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_3_rsci_douta_d,
      din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_4_rsci_douta_d, din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_5_rsci_douta_d, din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_6_rsci_douta_d,
      din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_7_rsci_douta_d, din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_8_rsci_douta_d, din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_9_rsci_douta_d,
      din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_10_rsci_douta_d, din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_11_rsci_douta_d, din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_12_rsci_douta_d,
      din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_13_rsci_douta_d, din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_14_rsci_douta_d, din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_15_rsci_douta_d,
      din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_16_rsci_douta_d, din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_17_rsci_douta_d, din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d, din_0_rsci_addra_d_pff
);
  input clk;
  input rst;
  input din_0_rsc_req_vz;
  output din_0_rsc_rls_lz;
  input din_1_rsc_req_vz;
  output din_1_rsc_rls_lz;
  input din_2_rsc_req_vz;
  output din_2_rsc_rls_lz;
  input din_3_rsc_req_vz;
  output din_3_rsc_rls_lz;
  input din_4_rsc_req_vz;
  output din_4_rsc_rls_lz;
  input din_5_rsc_req_vz;
  output din_5_rsc_rls_lz;
  input din_6_rsc_req_vz;
  output din_6_rsc_rls_lz;
  input din_7_rsc_req_vz;
  output din_7_rsc_rls_lz;
  input din_8_rsc_req_vz;
  output din_8_rsc_rls_lz;
  input din_9_rsc_req_vz;
  output din_9_rsc_rls_lz;
  input din_10_rsc_req_vz;
  output din_10_rsc_rls_lz;
  input din_11_rsc_req_vz;
  output din_11_rsc_rls_lz;
  input din_12_rsc_req_vz;
  output din_12_rsc_rls_lz;
  input din_13_rsc_req_vz;
  output din_13_rsc_rls_lz;
  input din_14_rsc_req_vz;
  output din_14_rsc_rls_lz;
  input din_15_rsc_req_vz;
  output din_15_rsc_rls_lz;
  input din_16_rsc_req_vz;
  output din_16_rsc_rls_lz;
  input din_17_rsc_req_vz;
  output din_17_rsc_rls_lz;
  output [511:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;
  input [63:0] din_0_rsci_douta_d;
  output din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_1_rsci_douta_d;
  output din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_2_rsci_douta_d;
  output din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_3_rsci_douta_d;
  output din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_4_rsci_douta_d;
  output din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_5_rsci_douta_d;
  output din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_6_rsci_douta_d;
  output din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_7_rsci_douta_d;
  output din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_8_rsci_douta_d;
  output din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_9_rsci_douta_d;
  output din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_10_rsci_douta_d;
  output din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_11_rsci_douta_d;
  output din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_12_rsci_douta_d;
  output din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_13_rsci_douta_d;
  output din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_14_rsci_douta_d;
  output din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_15_rsci_douta_d;
  output din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_16_rsci_douta_d;
  output din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] din_17_rsci_douta_d;
  output din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [6:0] din_0_rsci_addra_d_pff;
  wire [7:0] nl_din_0_rsci_addra_d_pff;


  // Interconnect Declarations
  wire core_wen;
  wire [15:0] din_0_rsci_douta_d_mxwt;
  wire core_wten;
  wire [15:0] din_1_rsci_douta_d_mxwt;
  wire [15:0] din_2_rsci_douta_d_mxwt;
  wire [15:0] din_3_rsci_douta_d_mxwt;
  wire [15:0] din_4_rsci_douta_d_mxwt;
  wire [15:0] din_5_rsci_douta_d_mxwt;
  wire [15:0] din_6_rsci_douta_d_mxwt;
  wire [15:0] din_7_rsci_douta_d_mxwt;
  wire [15:0] din_8_rsci_douta_d_mxwt;
  wire [15:0] din_9_rsci_douta_d_mxwt;
  wire [15:0] din_10_rsci_douta_d_mxwt;
  wire [15:0] din_11_rsci_douta_d_mxwt;
  wire [15:0] din_12_rsci_douta_d_mxwt;
  wire [15:0] din_13_rsci_douta_d_mxwt;
  wire [15:0] din_14_rsci_douta_d_mxwt;
  wire [15:0] din_15_rsci_douta_d_mxwt;
  wire [15:0] din_16_rsci_douta_d_mxwt;
  wire [15:0] din_17_rsci_douta_d_mxwt;
  wire dout_rsci_wen_comp;
  wire din_17_rsc_req_obj_wen_comp;
  wire din_16_rsc_req_obj_wen_comp;
  wire din_15_rsc_req_obj_wen_comp;
  wire din_14_rsc_req_obj_wen_comp;
  wire din_13_rsc_req_obj_wen_comp;
  wire din_12_rsc_req_obj_wen_comp;
  wire din_11_rsc_req_obj_wen_comp;
  wire din_10_rsc_req_obj_wen_comp;
  wire din_9_rsc_req_obj_wen_comp;
  wire din_8_rsc_req_obj_wen_comp;
  wire din_7_rsc_req_obj_wen_comp;
  wire din_6_rsc_req_obj_wen_comp;
  wire din_5_rsc_req_obj_wen_comp;
  wire din_4_rsc_req_obj_wen_comp;
  wire din_3_rsc_req_obj_wen_comp;
  wire din_2_rsc_req_obj_wen_comp;
  wire din_1_rsc_req_obj_wen_comp;
  wire din_0_rsc_req_obj_wen_comp;
  reg [15:0] dout_rsci_d_495_480;
  reg [15:0] dout_rsci_d_463_448;
  reg [15:0] dout_rsci_d_431_416;
  reg [15:0] dout_rsci_d_399_384;
  reg [15:0] dout_rsci_d_367_352;
  reg [15:0] dout_rsci_d_335_320;
  reg [15:0] dout_rsci_d_303_288;
  reg [15:0] dout_rsci_d_271_256;
  reg [15:0] dout_rsci_d_239_224;
  reg [15:0] dout_rsci_d_207_192;
  reg [15:0] dout_rsci_d_175_160;
  reg [15:0] dout_rsci_d_143_128;
  reg [15:0] dout_rsci_d_111_96;
  reg [15:0] dout_rsci_d_79_64;
  reg [15:0] dout_rsci_d_47_32;
  reg [15:0] dout_rsci_d_15_0;
  wire [1:0] fsm_output;
  wire [2:0] READ_for_acc_1_tmp;
  wire [3:0] nl_READ_for_acc_1_tmp;
  wire [6:0] READ_for_for_acc_1_tmp;
  wire [7:0] nl_READ_for_for_acc_1_tmp;
  wire or_dcpl_1;
  wire and_dcpl_9;
  reg exitL_exit_READ_sva;
  reg [1:0] READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_4;
  reg exit_READ_for_for_for_lpi_1_dfm_2;
  reg [1:0] READ_for_for_for_wy_idx_1_0_lpi_1_dfm_5;
  reg exit_READ_for_for_lpi_1_dfm_2;
  reg exit_READ_for_lpi_1_dfm_2;
  reg [1:0] READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_5;
  reg main_stage_0_2;
  reg [1:0] READ_for_k_idx_2_0_lpi_1_dfm_1_1_0_1;
  reg [5:0] READ_for_for_y_idx_6_0_lpi_1_dfm_3_5_0_1;
  wire READ_for_for_for_acc_tmp_2;
  wire READ_for_for_for_for_acc_tmp_2;
  wire exit_READ_for_for_lpi_1_dfm_2_mx0w0;
  wire lfst_exit_READ_for_for_1_lpi_1_dfm;
  wire lfst_exit_READ_lpi_1_dfm;
  wire [1:0] READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm;
  wire [1:0] READ_for_for_for_for_wx_idx_1_0_sva_1;
  wire [2:0] nl_READ_for_for_for_for_wx_idx_1_0_sva_1;
  reg reg_din_17_rsc_req_obj_oswt_cse;
  wire dout_and_cse;
  reg reg_din_17_rsc_rls_obj_ld_core_psct_cse;
  reg reg_dout_rsci_ld_core_psct_cse;
  reg reg_din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse;
  reg reg_din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse;
  reg reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse;
  wire READ_and_cse;
  wire nor_1_cse;
  wire or_7_cse;
  wire or_2_cse;
  wire din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire and_24_rmff;
  wire din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire and_18_rmff;
  wire din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire and_15_rmff;
  wire [5:0] READ_for_for_y_idx_6_0_lpi_1_dfm_5_0;
  wire [1:0] READ_for_for_for_wy_idx_1_0_lpi_1_dfm;
  wire [1:0] READ_for_for_for_acc_1_tmp;
  wire [2:0] nl_READ_for_for_for_acc_1_tmp;
  wire exit_READ_for_lpi_1_dfm_2_mx0w0;
  wire READ_for_for_for_for_else_unequal_tmp;
  wire READ_for_for_for_for_unequal_tmp;
  wire [1:0] READ_for_k_idx_2_0_lpi_1_dfm_1_0;
  wire READ_for_for_y_idx_and_2_cse;

  wire[0:0] READ_for_for_for_for_and_1_nl;
  wire[0:0] READ_for_for_for_for_not_9_nl;
  wire[0:0] READ_for_for_for_for_not_10_nl;
  wire[0:0] READ_for_for_for_for_not_8_nl;
  wire[0:0] READ_for_for_for_wy_idx_and_nl;
  wire[0:0] READ_for_for_y_idx_and_nl;
  wire[0:0] READ_for_for_READ_for_for_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [511:0] nl_READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_inst_dout_rsci_d;
  assign nl_READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_inst_dout_rsci_d =
      signext_512_496({dout_rsci_d_495_480 , ({{16{dout_rsci_d_463_448[15]}}, dout_rsci_d_463_448})
      , ({{16{dout_rsci_d_431_416[15]}}, dout_rsci_d_431_416}) , ({{16{dout_rsci_d_399_384[15]}},
      dout_rsci_d_399_384}) , ({{16{dout_rsci_d_367_352[15]}}, dout_rsci_d_367_352})
      , ({{16{dout_rsci_d_335_320[15]}}, dout_rsci_d_335_320}) , ({{16{dout_rsci_d_303_288[15]}},
      dout_rsci_d_303_288}) , ({{16{dout_rsci_d_271_256[15]}}, dout_rsci_d_271_256})
      , ({{16{dout_rsci_d_239_224[15]}}, dout_rsci_d_239_224}) , ({{16{dout_rsci_d_207_192[15]}},
      dout_rsci_d_207_192}) , ({{16{dout_rsci_d_175_160[15]}}, dout_rsci_d_175_160})
      , ({{16{dout_rsci_d_143_128[15]}}, dout_rsci_d_143_128}) , ({{16{dout_rsci_d_111_96[15]}},
      dout_rsci_d_111_96}) , ({{16{dout_rsci_d_79_64[15]}}, dout_rsci_d_79_64}) ,
      ({{16{dout_rsci_d_47_32[15]}}, dout_rsci_d_47_32}) , ({{16{dout_rsci_d_15_0[15]}},
      dout_rsci_d_15_0})});
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_0_rsci_douta_d(din_0_rsci_douta_d),
      .din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .din_0_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_0_rsci_douta_d_mxwt(din_0_rsci_douta_d_mxwt),
      .core_wten(core_wten),
      .din_0_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_1_rsci_douta_d(din_1_rsci_douta_d),
      .din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_1_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_1_rsci_douta_d_mxwt(din_1_rsci_douta_d_mxwt),
      .din_1_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_2_rsci_douta_d(din_2_rsci_douta_d),
      .din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_2_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_2_rsci_douta_d_mxwt(din_2_rsci_douta_d_mxwt),
      .din_2_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_3_rsci_douta_d(din_3_rsci_douta_d),
      .din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_3_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_3_rsci_douta_d_mxwt(din_3_rsci_douta_d_mxwt),
      .din_3_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_4_rsci_douta_d(din_4_rsci_douta_d),
      .din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_4_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_4_rsci_douta_d_mxwt(din_4_rsci_douta_d_mxwt),
      .din_4_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_5_rsci_douta_d(din_5_rsci_douta_d),
      .din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_5_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_5_rsci_douta_d_mxwt(din_5_rsci_douta_d_mxwt),
      .din_5_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_6_rsci_douta_d(din_6_rsci_douta_d),
      .din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_6_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_6_rsci_douta_d_mxwt(din_6_rsci_douta_d_mxwt),
      .din_6_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_7_rsci_douta_d(din_7_rsci_douta_d),
      .din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_7_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_7_rsci_douta_d_mxwt(din_7_rsci_douta_d_mxwt),
      .din_7_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_8_rsci_douta_d(din_8_rsci_douta_d),
      .din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_8_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_8_rsci_douta_d_mxwt(din_8_rsci_douta_d_mxwt),
      .din_8_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_9_rsci_douta_d(din_9_rsci_douta_d),
      .din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_9_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_9_rsci_douta_d_mxwt(din_9_rsci_douta_d_mxwt),
      .din_9_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_10_rsci_douta_d(din_10_rsci_douta_d),
      .din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_10_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_10_rsci_douta_d_mxwt(din_10_rsci_douta_d_mxwt),
      .din_10_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_11_rsci_douta_d(din_11_rsci_douta_d),
      .din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_11_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_11_rsci_douta_d_mxwt(din_11_rsci_douta_d_mxwt),
      .din_11_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_12_rsci_douta_d(din_12_rsci_douta_d),
      .din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_12_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_12_rsci_douta_d_mxwt(din_12_rsci_douta_d_mxwt),
      .din_12_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_13_rsci_douta_d(din_13_rsci_douta_d),
      .din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_13_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_13_rsci_douta_d_mxwt(din_13_rsci_douta_d_mxwt),
      .din_13_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_14_rsci_douta_d(din_14_rsci_douta_d),
      .din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_14_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_14_rsci_douta_d_mxwt(din_14_rsci_douta_d_mxwt),
      .din_14_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_15_rsci_douta_d(din_15_rsci_douta_d),
      .din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_15_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_15_rsci_douta_d_mxwt(din_15_rsci_douta_d_mxwt),
      .din_15_rsci_oswt_pff(and_24_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_16_rsci_douta_d(din_16_rsci_douta_d),
      .din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_16_rsci_oswt(reg_din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_16_rsci_douta_d_mxwt(din_16_rsci_douta_d_mxwt),
      .din_16_rsci_oswt_pff(and_18_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_17_rsci_douta_d(din_17_rsci_douta_d),
      .din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_17_rsci_oswt(reg_din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_17_rsci_douta_d_mxwt(din_17_rsci_douta_d_mxwt),
      .din_17_rsci_oswt_pff(and_15_rmff)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_rsc_z(dout_rsc_z),
      .dout_rsc_vz(dout_rsc_vz),
      .dout_rsc_lz(dout_rsc_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsci_oswt(reg_dout_rsci_ld_core_psct_cse),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_d(nl_READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_dout_rsci_inst_dout_rsci_d[511:0])
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_rls_obj_inst
      (
      .din_0_rsc_rls_lz(din_0_rsc_rls_lz),
      .core_wten(core_wten),
      .din_0_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_rls_obj_inst
      (
      .din_1_rsc_rls_lz(din_1_rsc_rls_lz),
      .core_wten(core_wten),
      .din_1_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_rls_obj_inst
      (
      .din_2_rsc_rls_lz(din_2_rsc_rls_lz),
      .core_wten(core_wten),
      .din_2_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_rls_obj_inst
      (
      .din_3_rsc_rls_lz(din_3_rsc_rls_lz),
      .core_wten(core_wten),
      .din_3_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_rls_obj_inst
      (
      .din_4_rsc_rls_lz(din_4_rsc_rls_lz),
      .core_wten(core_wten),
      .din_4_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_rls_obj_inst
      (
      .din_5_rsc_rls_lz(din_5_rsc_rls_lz),
      .core_wten(core_wten),
      .din_5_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_rls_obj_inst
      (
      .din_6_rsc_rls_lz(din_6_rsc_rls_lz),
      .core_wten(core_wten),
      .din_6_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_rls_obj_inst
      (
      .din_7_rsc_rls_lz(din_7_rsc_rls_lz),
      .core_wten(core_wten),
      .din_7_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_rls_obj_inst
      (
      .din_8_rsc_rls_lz(din_8_rsc_rls_lz),
      .core_wten(core_wten),
      .din_8_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_rls_obj_inst
      (
      .din_9_rsc_rls_lz(din_9_rsc_rls_lz),
      .core_wten(core_wten),
      .din_9_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_rls_obj_inst
      (
      .din_10_rsc_rls_lz(din_10_rsc_rls_lz),
      .core_wten(core_wten),
      .din_10_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_rls_obj_inst
      (
      .din_11_rsc_rls_lz(din_11_rsc_rls_lz),
      .core_wten(core_wten),
      .din_11_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_rls_obj_inst
      (
      .din_12_rsc_rls_lz(din_12_rsc_rls_lz),
      .core_wten(core_wten),
      .din_12_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_rls_obj_inst
      (
      .din_13_rsc_rls_lz(din_13_rsc_rls_lz),
      .core_wten(core_wten),
      .din_13_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_rls_obj_inst
      (
      .din_14_rsc_rls_lz(din_14_rsc_rls_lz),
      .core_wten(core_wten),
      .din_14_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_rls_obj_inst
      (
      .din_15_rsc_rls_lz(din_15_rsc_rls_lz),
      .core_wten(core_wten),
      .din_15_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_rls_obj_inst
      (
      .din_16_rsc_rls_lz(din_16_rsc_rls_lz),
      .core_wten(core_wten),
      .din_16_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_rls_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_rls_obj_inst
      (
      .din_17_rsc_rls_lz(din_17_rsc_rls_lz),
      .core_wten(core_wten),
      .din_17_rsc_rls_obj_iswt0(reg_din_17_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_17_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_17_rsc_req_vz(din_17_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_17_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_17_rsc_req_obj_wen_comp(din_17_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_16_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_16_rsc_req_vz(din_16_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_16_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_16_rsc_req_obj_wen_comp(din_16_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_15_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_15_rsc_req_vz(din_15_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_15_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_15_rsc_req_obj_wen_comp(din_15_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_14_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_14_rsc_req_vz(din_14_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_14_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_14_rsc_req_obj_wen_comp(din_14_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_13_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_13_rsc_req_vz(din_13_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_13_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_13_rsc_req_obj_wen_comp(din_13_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_12_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_12_rsc_req_vz(din_12_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_12_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_12_rsc_req_obj_wen_comp(din_12_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_11_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_11_rsc_req_vz(din_11_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_11_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_11_rsc_req_obj_wen_comp(din_11_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_10_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_10_rsc_req_vz(din_10_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_10_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_10_rsc_req_obj_wen_comp(din_10_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_9_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_9_rsc_req_vz(din_9_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_9_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_9_rsc_req_obj_wen_comp(din_9_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_8_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_8_rsc_req_vz(din_8_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_8_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_8_rsc_req_obj_wen_comp(din_8_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_7_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_7_rsc_req_vz(din_7_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_7_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_7_rsc_req_obj_wen_comp(din_7_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_6_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_6_rsc_req_vz(din_6_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_6_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_6_rsc_req_obj_wen_comp(din_6_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_5_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_5_rsc_req_vz(din_5_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_5_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_5_rsc_req_obj_wen_comp(din_5_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_4_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_4_rsc_req_vz(din_4_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_4_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_4_rsc_req_obj_wen_comp(din_4_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_3_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_3_rsc_req_vz(din_3_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_3_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_3_rsc_req_obj_wen_comp(din_3_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_2_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_2_rsc_req_vz(din_2_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_2_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_2_rsc_req_obj_wen_comp(din_2_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_1_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_1_rsc_req_vz(din_1_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_1_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_1_rsc_req_obj_wen_comp(din_1_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_din_0_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_0_rsc_req_vz(din_0_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_0_rsc_req_obj_oswt(reg_din_17_rsc_req_obj_oswt_cse),
      .din_0_rsc_req_obj_wen_comp(din_0_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_staller READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .din_17_rsc_req_obj_wen_comp(din_17_rsc_req_obj_wen_comp),
      .din_16_rsc_req_obj_wen_comp(din_16_rsc_req_obj_wen_comp),
      .din_15_rsc_req_obj_wen_comp(din_15_rsc_req_obj_wen_comp),
      .din_14_rsc_req_obj_wen_comp(din_14_rsc_req_obj_wen_comp),
      .din_13_rsc_req_obj_wen_comp(din_13_rsc_req_obj_wen_comp),
      .din_12_rsc_req_obj_wen_comp(din_12_rsc_req_obj_wen_comp),
      .din_11_rsc_req_obj_wen_comp(din_11_rsc_req_obj_wen_comp),
      .din_10_rsc_req_obj_wen_comp(din_10_rsc_req_obj_wen_comp),
      .din_9_rsc_req_obj_wen_comp(din_9_rsc_req_obj_wen_comp),
      .din_8_rsc_req_obj_wen_comp(din_8_rsc_req_obj_wen_comp),
      .din_7_rsc_req_obj_wen_comp(din_7_rsc_req_obj_wen_comp),
      .din_6_rsc_req_obj_wen_comp(din_6_rsc_req_obj_wen_comp),
      .din_5_rsc_req_obj_wen_comp(din_5_rsc_req_obj_wen_comp),
      .din_4_rsc_req_obj_wen_comp(din_4_rsc_req_obj_wen_comp),
      .din_3_rsc_req_obj_wen_comp(din_3_rsc_req_obj_wen_comp),
      .din_2_rsc_req_obj_wen_comp(din_2_rsc_req_obj_wen_comp),
      .din_1_rsc_req_obj_wen_comp(din_1_rsc_req_obj_wen_comp),
      .din_0_rsc_req_obj_wen_comp(din_0_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_core_fsm READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_core_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign or_7_cse = or_dcpl_1 | (~ (READ_for_for_acc_1_tmp[6])) | (~ (READ_for_acc_1_tmp[2]));
  assign dout_and_cse = core_wen & main_stage_0_2;
  assign and_15_rmff = and_dcpl_9 & (~ exitL_exit_READ_sva) & (READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_4[1]);
  assign and_18_rmff = and_dcpl_9 & (~ exitL_exit_READ_sva) & (READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_4==2'b01);
  assign and_24_rmff = (exit_READ_for_for_for_lpi_1_dfm_2 | exit_READ_for_for_lpi_1_dfm_2
      | exit_READ_for_lpi_1_dfm_2 | (~((READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_4!=2'b00)))
      | exitL_exit_READ_sva) & (fsm_output[1]);
  assign READ_and_cse = core_wen & (~ (fsm_output[0]));
  assign or_2_cse = or_dcpl_1 | (~ (READ_for_for_acc_1_tmp[6]));
  assign READ_for_for_y_idx_and_2_cse = core_wen & or_7_cse;
  assign nor_1_cse = ~(READ_for_for_for_for_acc_tmp_2 | READ_for_for_for_acc_tmp_2);
  assign exit_READ_for_lpi_1_dfm_2_mx0w0 = (READ_for_acc_1_tmp[2]) & exit_READ_for_for_lpi_1_dfm_2_mx0w0;
  assign READ_for_for_READ_for_for_and_1_nl = (~ exit_READ_for_for_for_lpi_1_dfm_2)
      & lfst_exit_READ_for_for_1_lpi_1_dfm;
  assign READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm = MUX_v_2_2_2(2'b00, READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_4,
      (READ_for_for_READ_for_for_and_1_nl));
  assign READ_for_for_for_acc_tmp_2 = (READ_for_for_for_acc_1_tmp[0]) ^ (READ_for_for_for_acc_1_tmp[1]);
  assign exit_READ_for_for_lpi_1_dfm_2_mx0w0 = (READ_for_for_acc_1_tmp[6]) & nor_1_cse;
  assign READ_for_for_for_for_else_unequal_tmp = ~((READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_5==2'b01));
  assign READ_for_for_for_for_unequal_tmp = (READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_5!=2'b00);
  assign nl_READ_for_acc_1_tmp = conv_u2u_2_3(READ_for_k_idx_2_0_lpi_1_dfm_1_0) +
      3'b1;
  assign READ_for_acc_1_tmp = nl_READ_for_acc_1_tmp[2:0];
  assign READ_for_k_idx_2_0_lpi_1_dfm_1_0 = MUX_v_2_2_2(2'b00, READ_for_k_idx_2_0_lpi_1_dfm_1_1_0_1,
      lfst_exit_READ_lpi_1_dfm);
  assign nl_READ_for_for_acc_1_tmp = conv_u2u_6_7(READ_for_for_y_idx_6_0_lpi_1_dfm_5_0)
      + 7'b1;
  assign READ_for_for_acc_1_tmp = nl_READ_for_for_acc_1_tmp[6:0];
  assign READ_for_for_y_idx_6_0_lpi_1_dfm_5_0 = MUX_v_6_2_2(6'b000000, READ_for_for_y_idx_6_0_lpi_1_dfm_3_5_0_1,
      lfst_exit_READ_lpi_1_dfm);
  assign nl_READ_for_for_for_acc_1_tmp = READ_for_for_for_wy_idx_1_0_lpi_1_dfm +
      2'b1;
  assign READ_for_for_for_acc_1_tmp = nl_READ_for_for_for_acc_1_tmp[1:0];
  assign READ_for_for_for_wy_idx_1_0_lpi_1_dfm = MUX_v_2_2_2(2'b00, READ_for_for_for_wy_idx_1_0_lpi_1_dfm_5,
      lfst_exit_READ_for_for_1_lpi_1_dfm);
  assign READ_for_for_for_for_acc_tmp_2 = (READ_for_for_for_for_wx_idx_1_0_sva_1[0])
      ^ (READ_for_for_for_for_wx_idx_1_0_sva_1[1]);
  assign nl_READ_for_for_for_for_wx_idx_1_0_sva_1 = READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm
      + 2'b1;
  assign READ_for_for_for_for_wx_idx_1_0_sva_1 = nl_READ_for_for_for_for_wx_idx_1_0_sva_1[1:0];
  assign lfst_exit_READ_for_for_1_lpi_1_dfm = (~ exit_READ_for_for_lpi_1_dfm_2) &
      lfst_exit_READ_lpi_1_dfm;
  assign lfst_exit_READ_lpi_1_dfm = ~(exit_READ_for_lpi_1_dfm_2 | exitL_exit_READ_sva);
  assign or_dcpl_1 = READ_for_for_for_for_acc_tmp_2 | READ_for_for_for_acc_tmp_2;
  assign and_dcpl_9 = ~(exit_READ_for_for_for_lpi_1_dfm_2 | exit_READ_for_for_lpi_1_dfm_2
      | exit_READ_for_lpi_1_dfm_2);
  assign nl_din_0_rsci_addra_d_pff = conv_u2u_6_7(READ_for_for_y_idx_6_0_lpi_1_dfm_5_0)
      + conv_u2u_2_7(READ_for_for_for_wy_idx_1_0_lpi_1_dfm);
  assign din_0_rsci_addra_d_pff = nl_din_0_rsci_addra_d_pff[6:0];
  assign din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      reg_din_17_rsc_req_obj_oswt_cse <= 1'b0;
      reg_din_17_rsc_rls_obj_ld_core_psct_cse <= 1'b0;
      reg_dout_rsci_ld_core_psct_cse <= 1'b0;
      reg_din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse <= 1'b0;
      reg_din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse <= 1'b0;
      reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse <= 1'b0;
      READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_5 <= 2'b0;
      main_stage_0_2 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_din_17_rsc_req_obj_oswt_cse <= ~(or_7_cse & (fsm_output[1]));
      reg_din_17_rsc_rls_obj_ld_core_psct_cse <= nor_1_cse & (READ_for_for_acc_1_tmp[6])
          & (READ_for_acc_1_tmp[2]) & (fsm_output[1]);
      reg_dout_rsci_ld_core_psct_cse <= main_stage_0_2;
      reg_din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse <= and_15_rmff;
      reg_din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse <= and_18_rmff;
      reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse <= and_24_rmff;
      READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_5 <= READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm;
      main_stage_0_2 <= fsm_output[1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_d_15_0 <= 16'b0;
      dout_rsci_d_47_32 <= 16'b0;
      dout_rsci_d_79_64 <= 16'b0;
      dout_rsci_d_111_96 <= 16'b0;
      dout_rsci_d_143_128 <= 16'b0;
      dout_rsci_d_175_160 <= 16'b0;
      dout_rsci_d_207_192 <= 16'b0;
      dout_rsci_d_239_224 <= 16'b0;
      dout_rsci_d_271_256 <= 16'b0;
      dout_rsci_d_303_288 <= 16'b0;
      dout_rsci_d_335_320 <= 16'b0;
      dout_rsci_d_367_352 <= 16'b0;
      dout_rsci_d_399_384 <= 16'b0;
      dout_rsci_d_431_416 <= 16'b0;
      dout_rsci_d_463_448 <= 16'b0;
      dout_rsci_d_495_480 <= 16'b0;
    end
    else if ( dout_and_cse ) begin
      dout_rsci_d_15_0 <= MUX1HOT_v_16_3_2(din_0_rsci_douta_d_mxwt, din_16_rsci_douta_d_mxwt,
          din_17_rsci_douta_d_mxwt, {(~ READ_for_for_for_for_unequal_tmp) , (~ READ_for_for_for_for_else_unequal_tmp)
          , (READ_for_for_for_for_and_1_nl)});
      dout_rsci_d_47_32 <= MUX_v_16_2_2(16'b0000000000000000, din_1_rsci_douta_d_mxwt,
          (READ_for_for_for_for_not_9_nl));
      dout_rsci_d_79_64 <= MUX_v_16_2_2(16'b0000000000000000, din_2_rsci_douta_d_mxwt,
          (READ_for_for_for_for_not_10_nl));
      dout_rsci_d_111_96 <= MUX_v_16_2_2(16'b0000000000000000, din_3_rsci_douta_d_mxwt,
          (READ_for_for_for_for_not_8_nl));
      dout_rsci_d_143_128 <= din_4_rsci_douta_d_mxwt;
      dout_rsci_d_175_160 <= din_5_rsci_douta_d_mxwt;
      dout_rsci_d_207_192 <= din_6_rsci_douta_d_mxwt;
      dout_rsci_d_239_224 <= din_7_rsci_douta_d_mxwt;
      dout_rsci_d_271_256 <= din_8_rsci_douta_d_mxwt;
      dout_rsci_d_303_288 <= din_9_rsci_douta_d_mxwt;
      dout_rsci_d_335_320 <= din_10_rsci_douta_d_mxwt;
      dout_rsci_d_367_352 <= din_11_rsci_douta_d_mxwt;
      dout_rsci_d_399_384 <= din_12_rsci_douta_d_mxwt;
      dout_rsci_d_431_416 <= din_13_rsci_douta_d_mxwt;
      dout_rsci_d_463_448 <= din_14_rsci_douta_d_mxwt;
      dout_rsci_d_495_480 <= din_15_rsci_douta_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exitL_exit_READ_sva <= 1'b1;
      exit_READ_for_lpi_1_dfm_2 <= 1'b0;
      exit_READ_for_for_lpi_1_dfm_2 <= 1'b0;
      exit_READ_for_for_for_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( READ_and_cse ) begin
      exitL_exit_READ_sva <= exit_READ_for_lpi_1_dfm_2_mx0w0;
      exit_READ_for_lpi_1_dfm_2 <= exit_READ_for_lpi_1_dfm_2_mx0w0;
      exit_READ_for_for_lpi_1_dfm_2 <= exit_READ_for_for_lpi_1_dfm_2_mx0w0;
      exit_READ_for_for_for_lpi_1_dfm_2 <= nor_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_4 <= 2'b0;
    end
    else if ( core_wen & or_dcpl_1 ) begin
      READ_for_for_for_for_wx_idx_1_0_lpi_1_dfm_4 <= MUX_v_2_2_2((signext_2_1(~ READ_for_for_for_acc_tmp_2)),
          READ_for_for_for_for_wx_idx_1_0_sva_1, READ_for_for_for_for_acc_tmp_2);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      READ_for_for_for_wy_idx_1_0_lpi_1_dfm_5 <= 2'b0;
    end
    else if ( core_wen & or_2_cse ) begin
      READ_for_for_for_wy_idx_1_0_lpi_1_dfm_5 <= MUX1HOT_v_2_3_2((signext_2_1(READ_for_for_acc_1_tmp[6])),
          READ_for_for_for_acc_1_tmp, READ_for_for_for_wy_idx_1_0_lpi_1_dfm, {(~
          or_dcpl_1) , (READ_for_for_for_wy_idx_and_nl) , READ_for_for_for_for_acc_tmp_2});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      READ_for_for_y_idx_6_0_lpi_1_dfm_3_5_0_1 <= 6'b0;
      READ_for_k_idx_2_0_lpi_1_dfm_1_1_0_1 <= 2'b0;
    end
    else if ( READ_for_for_y_idx_and_2_cse ) begin
      READ_for_for_y_idx_6_0_lpi_1_dfm_3_5_0_1 <= MUX1HOT_v_6_3_2((signext_6_1(READ_for_acc_1_tmp[2])),
          (READ_for_for_acc_1_tmp[5:0]), READ_for_for_y_idx_6_0_lpi_1_dfm_5_0, {(~
          or_2_cse) , (READ_for_for_y_idx_and_nl) , or_dcpl_1});
      READ_for_k_idx_2_0_lpi_1_dfm_1_1_0_1 <= MUX_v_2_2_2((READ_for_acc_1_tmp[1:0]),
          READ_for_k_idx_2_0_lpi_1_dfm_1_0, or_2_cse);
    end
  end
  assign READ_for_for_for_for_and_1_nl = READ_for_for_for_for_else_unequal_tmp &
      READ_for_for_for_for_unequal_tmp;
  assign READ_for_for_for_for_not_9_nl = ~ READ_for_for_for_for_unequal_tmp;
  assign READ_for_for_for_for_not_10_nl = ~ READ_for_for_for_for_unequal_tmp;
  assign READ_for_for_for_for_not_8_nl = ~ READ_for_for_for_for_unequal_tmp;
  assign READ_for_for_for_wy_idx_and_nl = (~ READ_for_for_for_for_acc_tmp_2) & or_dcpl_1;
  assign READ_for_for_y_idx_and_nl = (~ or_dcpl_1) & or_2_cse;

  function [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function [511:0] signext_512_496;
    input [495:0] vector;
  begin
    signext_512_496= {{16{vector[495]}}, vector};
  end
  endfunction


  function [5:0] signext_6_1;
    input [0:0] vector;
  begin
    signext_6_1= {{5{vector[0]}}, vector};
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function  [6:0] conv_u2u_2_7 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_7 = {{5{1'b0}}, vector};
  end
  endfunction


  function  [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, dout_rsc_req_vz, dout_rsc_rls_lz,
      dout_rsci_addra_d, dout_rsci_addrb_d, dout_rsci_dinb_d, dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d
);
  input clk;
  input rst;
  input [63:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  input dout_rsc_req_vz;
  output dout_rsc_rls_lz;
  output [6:0] dout_rsci_addra_d;
  output [6:0] dout_rsci_addrb_d;
  output [63:0] dout_rsci_dinb_d;
  output dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;


  // Interconnect Declarations
  wire core_wen;
  wire din_rsci_wen_comp;
  wire [63:0] din_rsci_d_mxwt;
  wire core_wten;
  wire dout_rsc_req_obj_wen_comp;
  wire [1:0] fsm_output;
  wire [2:0] for_acc_1_tmp;
  wire [3:0] nl_for_acc_1_tmp;
  reg exitL_exit_for_sva;
  reg [3:0] for_for_for_wx_idx_3_0_lpi_1_dfm_4;
  reg exit_for_lpi_1_dfm_2;
  reg [1:0] for_k_idx_2_0_lpi_1_dfm_1_1_0_1;
  reg reg_dout_rsc_req_obj_oswt_cse;
  reg reg_dout_rsc_rls_obj_ld_core_psct_cse;
  reg reg_din_rsci_ld_core_psct_cse;
  wire for_and_cse;
  wire or_1_cse;
  wire [6:0] dout_rsci_addra_d_reg;
  wire [2:0] for_for_for_acc_6_rmff;
  wire [3:0] nl_for_for_for_acc_6_rmff;
  wire [6:0] dout_rsci_addrb_d_reg;
  wire dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [3:0] for_for_for_acc_5_psp;
  wire [4:0] nl_for_for_for_acc_5_psp;
  wire exit_for_lpi_1_dfm_2_mx0w0;
  wire [1:0] for_k_idx_2_0_lpi_1_dfm_1_0;
  wire [3:0] for_for_for_wx_idx_3_0_sva_1;
  wire [4:0] nl_for_for_for_wx_idx_3_0_sva_1;
  wire [3:0] for_for_for_wx_idx_3_0_lpi_1_dfm;
  wire for_for_for_wx_idx_and_cse;
  wire for_for_for_acc_itm_3_1;

  wire[0:0] for_not_7_nl;
  wire[3:0] for_for_for_acc_nl;
  wire[4:0] nl_for_for_for_acc_nl;
  wire[0:0] nor_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [6:0] nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_dout_rsci_addra_d_core;
  assign nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_dout_rsci_addra_d_core
      = {1'b0 , for_for_for_acc_6_rmff , (for_for_for_acc_5_psp[2:0])};
  wire [6:0] nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_dout_rsci_addrb_d_core;
  assign nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_dout_rsci_addrb_d_core
      = {1'b0 , for_for_for_acc_6_rmff , (for_for_for_acc_5_psp[2:0])};
  wire [0:0] nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_dout_rsci_iswt0_pff;
  assign nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_dout_rsci_iswt0_pff
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_core_wten_pff;
  assign nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_core_wten_pff
      = ~ core_wen;
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_din_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(din_rsc_z),
      .din_rsc_vz(din_rsc_vz),
      .din_rsc_lz(din_rsc_lz),
      .core_wen(core_wen),
      .din_rsci_oswt(reg_din_rsci_ld_core_psct_cse),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_d_mxwt(din_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1 WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst
      (
      .dout_rsci_addra_d(dout_rsci_addra_d_reg),
      .dout_rsci_addrb_d(dout_rsci_addrb_d_reg),
      .dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .dout_rsci_addra_d_core(nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_dout_rsci_addra_d_core[6:0]),
      .dout_rsci_addrb_d_core(nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_dout_rsci_addrb_d_core[6:0]),
      .dout_rsci_iswt0_pff(nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_dout_rsci_iswt0_pff[0:0]),
      .core_wten_pff(nl_WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsci_1_inst_core_wten_pff[0:0])
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_rls_obj WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_rls_obj_inst
      (
      .dout_rsc_rls_lz(dout_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_rsc_rls_obj_iswt0(reg_dout_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_dout_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_rsc_req_vz(dout_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsc_req_obj_oswt(reg_dout_rsc_req_obj_oswt_cse),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_staller WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .core_wten(core_wten),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_core_fsm WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_core_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign nl_for_for_for_acc_6_rmff = conv_u2u_1_3(for_for_for_acc_5_psp[3]) + conv_u2u_2_3(for_k_idx_2_0_lpi_1_dfm_1_0);
  assign for_for_for_acc_6_rmff = nl_for_for_for_acc_6_rmff[2:0];
  assign for_and_cse = core_wen & (~ (fsm_output[0]));
  assign for_for_for_wx_idx_and_cse = core_wen & or_1_cse;
  assign or_1_cse = for_for_for_acc_itm_3_1 | (~ (for_acc_1_tmp[2]));
  assign exit_for_lpi_1_dfm_2_mx0w0 = (for_acc_1_tmp[2]) & (~ for_for_for_acc_itm_3_1);
  assign nl_for_acc_1_tmp = conv_u2u_2_3(for_k_idx_2_0_lpi_1_dfm_1_0) + 3'b1;
  assign for_acc_1_tmp = nl_for_acc_1_tmp[2:0];
  assign for_not_7_nl = ~ exitL_exit_for_sva;
  assign for_k_idx_2_0_lpi_1_dfm_1_0 = MUX_v_2_2_2(2'b00, for_k_idx_2_0_lpi_1_dfm_1_1_0_1,
      (for_not_7_nl));
  assign nl_for_for_for_acc_nl = for_for_for_wx_idx_3_0_sva_1 + 4'b111;
  assign for_for_for_acc_nl = nl_for_for_for_acc_nl[3:0];
  assign for_for_for_acc_itm_3_1 = readslicef_4_1_3((for_for_for_acc_nl));
  assign nl_for_for_for_wx_idx_3_0_sva_1 = for_for_for_wx_idx_3_0_lpi_1_dfm + 4'b1;
  assign for_for_for_wx_idx_3_0_sva_1 = nl_for_for_for_wx_idx_3_0_sva_1[3:0];
  assign nor_nl = ~(exit_for_lpi_1_dfm_2 | exitL_exit_for_sva);
  assign for_for_for_wx_idx_3_0_lpi_1_dfm = MUX_v_4_2_2(4'b0000, for_for_for_wx_idx_3_0_lpi_1_dfm_4,
      (nor_nl));
  assign nl_for_for_for_acc_5_psp = for_for_for_wx_idx_3_0_lpi_1_dfm + conv_u2u_2_4(for_k_idx_2_0_lpi_1_dfm_1_0);
  assign for_for_for_acc_5_psp = nl_for_for_for_acc_5_psp[3:0];
  assign dout_rsci_addra_d = dout_rsci_addra_d_reg;
  assign dout_rsci_addrb_d = dout_rsci_addrb_d_reg;
  assign dout_rsci_dinb_d = din_rsci_d_mxwt;
  assign dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      reg_dout_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_rsc_rls_obj_ld_core_psct_cse <= 1'b0;
      reg_din_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_dout_rsc_req_obj_oswt_cse <= ~(or_1_cse & (fsm_output[1]));
      reg_dout_rsc_rls_obj_ld_core_psct_cse <= (~ for_for_for_acc_itm_3_1) & (for_acc_1_tmp[2])
          & (fsm_output[1]);
      reg_din_rsci_ld_core_psct_cse <= 1'b1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exitL_exit_for_sva <= 1'b1;
      exit_for_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( for_and_cse ) begin
      exitL_exit_for_sva <= exit_for_lpi_1_dfm_2_mx0w0;
      exit_for_lpi_1_dfm_2 <= exit_for_lpi_1_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_wx_idx_3_0_lpi_1_dfm_4 <= 4'b0;
      for_k_idx_2_0_lpi_1_dfm_1_1_0_1 <= 2'b0;
    end
    else if ( for_for_for_wx_idx_and_cse ) begin
      for_for_for_wx_idx_3_0_lpi_1_dfm_4 <= MUX_v_4_2_2((signext_4_1(for_acc_1_tmp[2])),
          for_for_for_wx_idx_3_0_sva_1, for_for_for_acc_itm_3_1);
      for_k_idx_2_0_lpi_1_dfm_1_1_0_1 <= MUX_v_2_2_2((for_acc_1_tmp[1:0]), for_k_idx_2_0_lpi_1_dfm_1_0,
          for_for_for_acc_itm_3_1);
    end
  end

  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function [3:0] signext_4_1;
    input [0:0] vector;
  begin
    signext_4_1= {{3{vector[0]}}, vector};
  end
  endfunction


  function  [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function  [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core (
  clk, rst, din_rsc_req_vz, din_rsc_rls_lz, dout_rsc_z, dout_rsc_vz, dout_rsc_lz,
      din_rsci_addra_d, din_rsci_addrb_d, din_rsci_douta_d, din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d
);
  input clk;
  input rst;
  input din_rsc_req_vz;
  output din_rsc_rls_lz;
  output [63:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;
  output [6:0] din_rsci_addra_d;
  output [6:0] din_rsci_addrb_d;
  input [63:0] din_rsci_douta_d;
  output din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations
  wire core_wen;
  wire [63:0] din_rsci_douta_d_mxwt;
  wire core_wten;
  wire dout_rsci_wen_comp;
  reg [63:0] dout_rsci_d;
  wire din_rsc_req_obj_wen_comp;
  wire [1:0] fsm_output;
  wire [2:0] for_acc_1_tmp;
  wire [3:0] nl_for_acc_1_tmp;
  reg exitL_exit_for_sva;
  reg [3:0] READ_for_wx_idx_3_0_lpi_1_dfm_4;
  reg exit_for_lpi_1_dfm_2;
  reg [1:0] for_k_idx_2_0_lpi_1_dfm_1_1_0_1;
  reg reg_din_rsc_req_obj_oswt_cse;
  reg reg_din_rsc_rls_obj_ld_core_psct_cse;
  reg reg_dout_rsci_ld_core_psct_cse;
  reg reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse;
  wire for_and_cse;
  wire or_1_cse;
  wire [6:0] din_rsci_addra_d_reg;
  wire [2:0] READ_for_acc_8_rmff;
  wire [3:0] nl_READ_for_acc_8_rmff;
  wire [6:0] din_rsci_addrb_d_reg;
  wire din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire [3:0] READ_for_acc_7_psp;
  wire [4:0] nl_READ_for_acc_7_psp;
  wire exit_for_lpi_1_dfm_2_mx0w0;
  wire [1:0] for_k_idx_2_0_lpi_1_dfm_1_0;
  wire [3:0] READ_for_wx_idx_3_0_sva_1;
  wire [4:0] nl_READ_for_wx_idx_3_0_sva_1;
  wire [3:0] READ_for_wx_idx_3_0_lpi_1_dfm;
  wire READ_for_wx_idx_and_cse;
  wire READ_for_acc_itm_3_1;

  wire[0:0] for_not_7_nl;
  wire[3:0] READ_for_acc_nl;
  wire[4:0] nl_READ_for_acc_nl;
  wire[0:0] nor_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [6:0] nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_inst_din_rsci_addra_d_core;
  assign nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_inst_din_rsci_addra_d_core
      = {1'b0 , READ_for_acc_8_rmff , (READ_for_acc_7_psp[2:0])};
  wire [6:0] nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_inst_din_rsci_addrb_d_core;
  assign nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_inst_din_rsci_addrb_d_core
      = {1'b0 , READ_for_acc_8_rmff , (READ_for_acc_7_psp[2:0])};
  wire [0:0] nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_inst_din_rsci_oswt_pff;
  assign nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_inst_din_rsci_oswt_pff
      = fsm_output[1];
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1 READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsci_addra_d(din_rsci_addra_d_reg),
      .din_rsci_addrb_d(din_rsci_addrb_d_reg),
      .din_rsci_douta_d(din_rsci_douta_d),
      .din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .din_rsci_oswt(reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_rsci_addra_d_core(nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_inst_din_rsci_addra_d_core[6:0]),
      .din_rsci_addrb_d_core(nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_inst_din_rsci_addrb_d_core[6:0]),
      .din_rsci_douta_d_mxwt(din_rsci_douta_d_mxwt),
      .core_wten(core_wten),
      .din_rsci_oswt_pff(nl_READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsci_1_inst_din_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_dout_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_rsc_z(dout_rsc_z),
      .dout_rsc_vz(dout_rsc_vz),
      .dout_rsc_lz(dout_rsc_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsci_oswt(reg_dout_rsci_ld_core_psct_cse),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_d(dout_rsci_d)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_rls_obj READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_rls_obj_inst
      (
      .din_rsc_rls_lz(din_rsc_rls_lz),
      .core_wten(core_wten),
      .din_rsc_rls_obj_iswt0(reg_din_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_din_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_req_vz(din_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_rsc_req_obj_oswt(reg_din_rsc_req_obj_oswt_cse),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_staller READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_core_fsm READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_core_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign nl_READ_for_acc_8_rmff = conv_u2u_1_3(READ_for_acc_7_psp[3]) + conv_u2u_2_3(for_k_idx_2_0_lpi_1_dfm_1_0);
  assign READ_for_acc_8_rmff = nl_READ_for_acc_8_rmff[2:0];
  assign for_and_cse = core_wen & (~ (fsm_output[0]));
  assign READ_for_wx_idx_and_cse = core_wen & or_1_cse;
  assign or_1_cse = READ_for_acc_itm_3_1 | (~ (for_acc_1_tmp[2]));
  assign exit_for_lpi_1_dfm_2_mx0w0 = (for_acc_1_tmp[2]) & (~ READ_for_acc_itm_3_1);
  assign nl_for_acc_1_tmp = conv_u2u_2_3(for_k_idx_2_0_lpi_1_dfm_1_0) + 3'b1;
  assign for_acc_1_tmp = nl_for_acc_1_tmp[2:0];
  assign for_not_7_nl = ~ exitL_exit_for_sva;
  assign for_k_idx_2_0_lpi_1_dfm_1_0 = MUX_v_2_2_2(2'b00, for_k_idx_2_0_lpi_1_dfm_1_1_0_1,
      (for_not_7_nl));
  assign nl_READ_for_acc_nl = READ_for_wx_idx_3_0_sva_1 + 4'b111;
  assign READ_for_acc_nl = nl_READ_for_acc_nl[3:0];
  assign READ_for_acc_itm_3_1 = readslicef_4_1_3((READ_for_acc_nl));
  assign nl_READ_for_wx_idx_3_0_sva_1 = READ_for_wx_idx_3_0_lpi_1_dfm + 4'b1;
  assign READ_for_wx_idx_3_0_sva_1 = nl_READ_for_wx_idx_3_0_sva_1[3:0];
  assign nor_nl = ~(exit_for_lpi_1_dfm_2 | exitL_exit_for_sva);
  assign READ_for_wx_idx_3_0_lpi_1_dfm = MUX_v_4_2_2(4'b0000, READ_for_wx_idx_3_0_lpi_1_dfm_4,
      (nor_nl));
  assign nl_READ_for_acc_7_psp = READ_for_wx_idx_3_0_lpi_1_dfm + conv_u2u_2_4(for_k_idx_2_0_lpi_1_dfm_1_0);
  assign READ_for_acc_7_psp = nl_READ_for_acc_7_psp[3:0];
  assign din_rsci_addra_d = din_rsci_addra_d_reg;
  assign din_rsci_addrb_d = din_rsci_addrb_d_reg;
  assign din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      reg_din_rsc_req_obj_oswt_cse <= 1'b0;
      reg_din_rsc_rls_obj_ld_core_psct_cse <= 1'b0;
      reg_dout_rsci_ld_core_psct_cse <= 1'b0;
      reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_din_rsc_req_obj_oswt_cse <= ~(or_1_cse & (fsm_output[1]));
      reg_din_rsc_rls_obj_ld_core_psct_cse <= (~ READ_for_acc_itm_3_1) & (for_acc_1_tmp[2])
          & (fsm_output[1]);
      reg_dout_rsci_ld_core_psct_cse <= reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse;
      reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse <= fsm_output[1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_d <= 64'b0;
    end
    else if ( core_wen & reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse
        ) begin
      dout_rsci_d <= din_rsci_douta_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exitL_exit_for_sva <= 1'b1;
      exit_for_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( for_and_cse ) begin
      exitL_exit_for_sva <= exit_for_lpi_1_dfm_2_mx0w0;
      exit_for_lpi_1_dfm_2 <= exit_for_lpi_1_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      READ_for_wx_idx_3_0_lpi_1_dfm_4 <= 4'b0;
      for_k_idx_2_0_lpi_1_dfm_1_1_0_1 <= 2'b0;
    end
    else if ( READ_for_wx_idx_and_cse ) begin
      READ_for_wx_idx_3_0_lpi_1_dfm_4 <= MUX_v_4_2_2((signext_4_1(for_acc_1_tmp[2])),
          READ_for_wx_idx_3_0_sva_1, READ_for_acc_itm_3_1);
      for_k_idx_2_0_lpi_1_dfm_1_1_0_1 <= MUX_v_2_2_2((for_acc_1_tmp[1:0]), for_k_idx_2_0_lpi_1_dfm_1_0,
          READ_for_acc_itm_3_1);
    end
  end

  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function [3:0] signext_4_1;
    input [0:0] vector;
  begin
    signext_4_1= {{3{vector[0]}}, vector};
  end
  endfunction


  function  [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function  [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array_core
// ------------------------------------------------------------------


module systolic_array_core (
  clk, rst, input_rsc_z, input_rsc_vz, input_rsc_lz, weight_rsc_z, weight_rsc_vz,
      weight_rsc_lz, output_rsc_z, output_rsc_vz, output_rsc_lz
);
  input clk;
  input rst;
  input [511:0] input_rsc_z;
  input input_rsc_vz;
  output input_rsc_lz;
  input [63:0] weight_rsc_z;
  input weight_rsc_vz;
  output weight_rsc_lz;
  output [1023:0] output_rsc_z;
  input output_rsc_vz;
  output output_rsc_lz;


  // Interconnect Declarations
  wire core_wen;
  wire input_rsci_wen_comp;
  wire [255:0] input_rsci_d_mxwt;
  wire core_wten;
  wire weight_rsci_wen_comp;
  wire [31:0] weight_rsci_d_mxwt;
  wire output_rsci_wen_comp;
  reg [1023:0] output_rsci_d;
  wire [1:0] WY_mux_6_tmp;
  wire COMP_and_13_tmp;
  wire [6:0] for_for_acc_1_tmp;
  wire [7:0] nl_for_for_acc_1_tmp;
  wire [4:0] for_for_for_1_acc_1_tmp;
  wire [5:0] nl_for_for_for_1_acc_1_tmp;
  wire for_for_for_1_nand_2_tmp;
  wire [2:0] for_acc_2_tmp;
  wire [3:0] nl_for_acc_2_tmp;
  wire [1:0] for_for_for_1_for_for_for_1_for_for_for_1_mux1h_1_tmp;
  wire and_dcpl_1;
  wire or_dcpl;
  wire or_tmp_4;
  wire or_tmp_5;
  wire mux_tmp;
  wire or_dcpl_7;
  wire or_dcpl_9;
  wire or_dcpl_13;
  wire or_dcpl_14;
  wire or_dcpl_15;
  wire and_dcpl_15;
  wire and_dcpl_27;
  wire or_dcpl_18;
  wire and_dcpl_36;
  wire or_tmp_16;
  wire and_tmp_2;
  wire or_tmp_19;
  wire and_dcpl_38;
  wire and_dcpl_48;
  wire or_dcpl_28;
  wire and_dcpl_59;
  wire or_dcpl_35;
  wire and_dcpl_61;
  wire and_dcpl_63;
  wire or_dcpl_38;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_68;
  wire and_dcpl_69;
  wire and_dcpl_70;
  wire and_dcpl_71;
  wire and_dcpl_72;
  wire and_dcpl_73;
  wire and_dcpl_74;
  wire and_dcpl_75;
  wire and_dcpl_76;
  wire and_dcpl_77;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_80;
  wire and_dcpl_81;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_87;
  wire and_dcpl_88;
  wire and_dcpl_89;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_92;
  wire and_dcpl_93;
  wire and_dcpl_94;
  wire and_dcpl_95;
  wire and_dcpl_96;
  wire and_dcpl_97;
  wire and_dcpl_98;
  wire and_dcpl_99;
  wire and_dcpl_100;
  wire and_dcpl_101;
  wire or_dcpl_50;
  wire or_dcpl_51;
  wire or_dcpl_70;
  wire or_dcpl_72;
  wire or_dcpl_76;
  reg [15:0] in_tmp_8_lpi_2;
  reg [15:0] in_tmp_7_lpi_2;
  reg [15:0] in_tmp_9_lpi_2;
  reg [15:0] in_tmp_6_lpi_2;
  reg [15:0] in_tmp_10_lpi_2;
  reg [15:0] in_tmp_5_lpi_2;
  reg [15:0] in_tmp_11_lpi_2;
  reg [15:0] in_tmp_4_lpi_2;
  reg [15:0] in_tmp_12_lpi_2;
  reg [15:0] in_tmp_3_lpi_2;
  reg [15:0] in_tmp_13_lpi_2;
  reg [15:0] in_tmp_2_lpi_2;
  reg [15:0] in_tmp_14_lpi_2;
  reg [15:0] in_tmp_1_lpi_2;
  reg [15:0] in_tmp_15_lpi_2;
  reg [15:0] weight_buf_value_1_1_15_0_lpi_1;
  reg [15:0] weight_buf_value_1_1_47_32_lpi_1;
  reg [15:0] weight_buf_value_1_0_15_0_lpi_1;
  reg [15:0] weight_buf_value_1_0_47_32_lpi_1;
  reg [15:0] weight_buf_value_1_2_15_0_lpi_1;
  reg [15:0] weight_buf_value_1_2_47_32_lpi_1;
  reg [15:0] weight_buf_value_0_2_15_0_lpi_1;
  reg [15:0] weight_buf_value_0_2_47_32_lpi_1;
  reg [15:0] weight_buf_value_2_0_15_0_lpi_1;
  reg [15:0] weight_buf_value_2_0_47_32_lpi_1;
  reg [15:0] weight_buf_value_0_1_15_0_lpi_1;
  reg [15:0] weight_buf_value_0_1_47_32_lpi_1;
  reg [15:0] weight_buf_value_2_1_15_0_lpi_1;
  reg [15:0] weight_buf_value_2_1_47_32_lpi_1;
  reg [15:0] weight_buf_value_0_0_15_0_lpi_1;
  reg [15:0] weight_buf_value_0_0_47_32_lpi_1;
  reg [15:0] weight_buf_value_2_2_15_0_lpi_1;
  reg [15:0] weight_buf_value_2_2_47_32_lpi_1;
  reg [6:0] for_for_row_6_0_lpi_3;
  reg lfst_exit_for_for_1_lpi_2;
  reg [31:0] out_tmp_value_0_31_0_lpi_2;
  reg [1:0] WY_wy_1_0_lpi_3;
  reg [1:0] WX_wx_1_0_lpi_3;
  reg lfst_exit_WX_1_lpi_1;
  reg exitL_exit_COL_1_COMP_lpi_1;
  reg [15:0] in_tmp_16_lpi_2;
  reg [15:0] pe_x_reg_0_lpi_2;
  reg COMP_i_0_1_lpi_1;
  reg [15:0] pe_x_reg_1_lpi_2;
  reg COMP_i_0_2_lpi_1;
  reg [15:0] pe_x_reg_2_lpi_2;
  reg COMP_i_0_3_lpi_1;
  reg [15:0] pe_x_reg_3_lpi_2;
  reg COMP_i_0_4_lpi_1;
  reg [15:0] pe_x_reg_4_lpi_2;
  reg COMP_i_0_5_lpi_1;
  reg [15:0] pe_x_reg_5_lpi_2;
  reg COMP_i_0_6_lpi_1;
  reg [15:0] pe_x_reg_6_lpi_2;
  reg COMP_i_0_7_lpi_1;
  reg [15:0] pe_x_reg_7_lpi_2;
  reg COMP_i_0_8_lpi_1;
  reg [15:0] pe_x_reg_8_lpi_2;
  reg COMP_i_0_9_lpi_1;
  reg [15:0] pe_x_reg_9_lpi_2;
  reg COMP_i_0_10_lpi_1;
  reg [15:0] pe_x_reg_10_lpi_2;
  reg COMP_i_0_11_lpi_1;
  reg [15:0] pe_x_reg_11_lpi_2;
  reg COMP_i_0_12_lpi_1;
  reg [15:0] pe_x_reg_12_lpi_2;
  reg COMP_i_0_13_lpi_1;
  reg [15:0] pe_x_reg_13_lpi_2;
  reg COMP_i_0_14_lpi_1;
  reg COMP_i_0_15_lpi_1;
  reg [31:0] pe_y_reg_value_7_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_7_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_8_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_8_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_6_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_6_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_9_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_9_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_5_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_5_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_10_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_10_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_4_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_4_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_11_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_11_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_3_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_3_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_12_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_12_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_2_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_2_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_13_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_13_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_1_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_1_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_14_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_14_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_0_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_0_63_32_lpi_2;
  reg [31:0] pe_y_reg_value_15_31_0_lpi_2;
  reg [31:0] pe_y_reg_value_15_63_32_lpi_2;
  reg COMP_i_0_lpi_1;
  reg for_for_for_1_for_q_0_lpi_2;
  reg exitL_exit_for_sva;
  reg WX_if_1_and_stg_1_0_sva;
  reg WX_if_1_and_stg_2_0_sva;
  reg WX_if_1_and_stg_1_3_sva;
  reg WX_if_1_and_stg_1_2_sva;
  reg WX_if_1_and_stg_1_1_sva;
  reg exit_WY_sva_2;
  reg exit_for_lpi_1_dfm_4;
  reg WX_and_1_psp_1;
  reg WX_and_3_psp_1;
  reg WX_and_5_psp_1;
  reg WX_and_7_psp_1;
  reg WX_and_9_psp_1;
  reg WX_and_11_psp_1;
  reg WX_and_13_psp_1;
  reg WX_and_15_psp_1;
  reg WX_and_17_psp_1;
  reg COMP_and_13_mdf_sva_5;
  reg COMP_and_13_mdf_sva_6;
  reg COMP_and_13_mdf_sva_7;
  reg WX_unequal_tmp_5;
  reg unequal_tmp_5;
  reg unequal_tmp_6;
  reg unequal_tmp_7;
  reg [31:0] out_tmp_value_15_31_0_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_15_63_32_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_14_31_0_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_14_63_32_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_13_31_0_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_13_63_32_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_12_31_0_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_12_63_32_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_11_31_0_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_11_63_32_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_10_31_0_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_10_63_32_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_9_31_0_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_9_63_32_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_8_31_0_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_8_63_32_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_7_31_0_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_7_63_32_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_6_31_0_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_6_63_32_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_5_31_0_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_5_63_32_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_4_31_0_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_4_63_32_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_3_31_0_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_3_63_32_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_2_31_0_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_2_63_32_lpi_1_dfm_12;
  reg [31:0] out_tmp_value_1_31_0_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_1_63_32_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_0_63_32_lpi_1_dfm_10;
  reg COMP_i_0_15_lpi_1_dfm_5;
  reg COMP_i_0_15_lpi_1_dfm_6;
  reg COMP_i_0_14_lpi_1_dfm_5;
  reg COMP_i_0_14_lpi_1_dfm_6;
  reg COMP_i_0_13_lpi_1_dfm_5;
  reg COMP_i_0_13_lpi_1_dfm_6;
  reg COMP_i_0_12_lpi_1_dfm_5;
  reg COMP_i_0_12_lpi_1_dfm_6;
  reg COMP_i_0_11_lpi_1_dfm_5;
  reg COMP_i_0_11_lpi_1_dfm_6;
  reg COMP_i_0_10_lpi_1_dfm_5;
  reg COMP_i_0_10_lpi_1_dfm_6;
  reg COMP_i_0_9_lpi_1_dfm_5;
  reg COMP_i_0_9_lpi_1_dfm_6;
  reg COMP_i_0_8_lpi_1_dfm_5;
  reg COMP_i_0_8_lpi_1_dfm_6;
  reg COMP_i_0_7_lpi_1_dfm_5;
  reg COMP_i_0_7_lpi_1_dfm_6;
  reg COMP_i_0_6_lpi_1_dfm_5;
  reg COMP_i_0_6_lpi_1_dfm_6;
  reg COMP_i_0_5_lpi_1_dfm_5;
  reg COMP_i_0_5_lpi_1_dfm_6;
  reg COMP_i_0_4_lpi_1_dfm_5;
  reg COMP_i_0_4_lpi_1_dfm_6;
  reg COMP_i_0_3_lpi_1_dfm_5;
  reg COMP_i_0_3_lpi_1_dfm_6;
  reg COMP_i_0_2_lpi_1_dfm_5;
  reg COMP_i_0_2_lpi_1_dfm_6;
  reg COMP_i_0_1_lpi_1_dfm_5;
  reg COMP_i_0_1_lpi_1_dfm_6;
  reg COMP_i_0_lpi_1_dfm_5;
  reg COMP_i_0_lpi_1_dfm_6;
  reg [15:0] in_tmp_16_lpi_1_dfm_5;
  reg [15:0] pe_x_reg_0_lpi_1_dfm_4;
  reg [6:0] for_for_row_6_0_lpi_1_dfm_9;
  reg lfst_exit_for_for_1_lpi_1_dfm_1;
  reg lfst_exit_for_for_1_lpi_1_dfm_4;
  reg [31:0] out_tmp_value_0_63_32_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_0_31_0_lpi_1_dfm_10;
  reg [31:0] out_tmp_value_1_63_32_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_1_31_0_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_2_63_32_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_2_31_0_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_3_63_32_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_3_31_0_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_4_63_32_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_4_31_0_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_5_63_32_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_5_31_0_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_6_63_32_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_6_31_0_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_7_63_32_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_7_31_0_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_8_63_32_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_8_31_0_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_9_63_32_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_9_31_0_lpi_1_dfm_13;
  reg [31:0] out_tmp_value_10_63_32_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_10_31_0_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_11_63_32_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_11_31_0_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_12_63_32_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_12_31_0_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_13_63_32_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_13_31_0_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_14_63_32_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_14_31_0_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_15_63_32_lpi_1_dfm_11;
  reg [31:0] out_tmp_value_15_31_0_lpi_1_dfm_11;
  reg for_for_for_1_equal_tmp_2;
  reg for_for_for_1_equal_tmp_10;
  reg for_for_for_1_equal_tmp_11;
  reg for_for_for_1_equal_tmp_5;
  reg for_for_for_1_equal_tmp_12;
  reg for_for_for_1_equal_tmp_13;
  reg exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  reg [15:0] COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000;
  reg for_for_for_1_nor_dfs_5;
  reg for_for_for_1_nor_dfs_6;
  reg for_for_for_1_nor_dfs_7;
  reg [15:0] mux_36_itm_2;
  reg [15:0] mux_37_itm_2;
  reg [15:0] mux_38_itm_2;
  reg [15:0] mux_39_itm_2;
  reg [15:0] mux_40_itm_2;
  reg [15:0] mux_41_itm_2;
  reg [15:0] mux_42_itm_2;
  reg [15:0] mux_43_itm_2;
  reg [15:0] mux_44_itm_2;
  reg [15:0] mux_45_itm_2;
  reg [15:0] mux_46_itm_2;
  reg [15:0] mux_47_itm_2;
  reg [15:0] mux_48_itm_2;
  reg [15:0] mux_63_itm_2;
  reg [31:0] COMP_mux_2_itm_2;
  reg [31:0] COMP_mux_3_itm_2;
  reg [31:0] COMP_mux_4_itm_2;
  reg [31:0] COMP_mux_5_itm_2;
  reg [31:0] COMP_mux_6_itm_2;
  reg [31:0] COMP_mux_7_itm_2;
  reg [31:0] COMP_mux_8_itm_2;
  reg [31:0] COMP_mux_9_itm_2;
  reg [31:0] COMP_mux_10_itm_2;
  reg [31:0] COMP_mux_11_itm_2;
  reg [31:0] COMP_mux_12_itm_2;
  reg [31:0] COMP_mux_13_itm_2;
  reg [31:0] COMP_mux_14_itm_2;
  reg [31:0] COMP_mux_15_itm_2;
  reg [31:0] COMP_mux_16_itm_2;
  reg [31:0] COMP_mux_17_itm_2;
  reg [31:0] COMP_mux_18_itm_2;
  reg [31:0] COMP_mux_19_itm_2;
  reg [31:0] COMP_mux_20_itm_2;
  reg [31:0] COMP_mux_21_itm_2;
  reg [31:0] COMP_mux_22_itm_2;
  reg [31:0] COMP_mux_23_itm_2;
  reg [31:0] COMP_mux_24_itm_2;
  reg [31:0] COMP_mux_25_itm_2;
  reg [31:0] COMP_mux_26_itm_2;
  reg [31:0] COMP_mux_27_itm_2;
  reg [31:0] COMP_mux_28_itm_2;
  reg [31:0] COMP_mux_29_itm_2;
  reg [31:0] COMP_mux_30_itm_2;
  reg [31:0] COMP_mux_31_itm_2;
  reg [31:0] COMP_mux_32_itm_2;
  reg [31:0] COMP_mux_33_itm_2;
  reg [1023:0] for_for_for_1_asn_itm_2;
  reg [5:0] for_for_row_slc_for_for_row_6_0_5_0_1_itm_3;
  reg [1:0] lfst_exit_for_for_for_1_lpi_1_dfm_1_st_4;
  reg [1:0] lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5;
  reg exit_for_for_for_1_lpi_1_dfm_1_st_3;
  reg exit_for_for_for_1_lpi_1_dfm_1_st_4;
  reg slc_lfst_exit_for_for_for_1_1_1_itm_4;
  reg main_stage_0_2;
  reg main_stage_0_3;
  reg main_stage_0_4;
  reg [1:0] for_ko_2_0_lpi_1_1_0_1;
  reg [3:0] for_for_for_1_k_4_0_lpi_1_3_0_1;
  reg lfst_exit_for_for_for_1_lpi_1_dfm_9_1_1;
  reg lfst_exit_for_for_for_1_lpi_1_dfm_10_1_1;
  reg for_for_row_6_0_lpi_1_dfm_6_6_1;
  reg for_for_row_6_0_lpi_1_dfm_7_6_1;
  reg PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_lo_conc_1_itm_2_5_1;
  reg out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1;
  reg lfst_exit_for_for_for_1_lpi_1_1_1;
  reg lfst_exit_for_for_for_1_lpi_1_0_1;
  reg [2:0] pref_pref_pref_6_3_0_1_lpi_1_3_1_1;
  reg pref_pref_pref_6_3_0_1_lpi_1_0_1;
  reg [2:0] WX_if_1_acc_decb_sva_3_1;
  reg [2:0] WX_if_1_acc_decb_sva_1_3_1_1;
  reg lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1;
  reg lfst_exit_for_for_for_1_lpi_1_dfm_st_1_0;
  reg lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1;
  reg lfst_exit_for_for_for_1_lpi_1_dfm_st_2_0_1;
  wire exit_WX_lpi_1_dfm_1;
  wire WY_unequal_tmp;
  wire lfst_exit_for_for_for_1_lpi_1_dfm_1;
  wire lfst_exit_for_for_for_1_lpi_1_dfm_0;
  wire exit_for_for_for_1_lpi_1_dfm_1;
  wire lfst_exit_for_for_1_lpi_1_dfm;
  wire lfst_exit_for_lpi_1_dfm;
  wire for_for_for_1_and_3_cse;
  wire for_for_for_1_and_4_m1c;
  wire for_for_for_1_and_96_cse;
  wire for_for_for_1_equal_tmp_1;
  wire for_for_for_1_and_95_cse;
  wire for_for_for_1_equal_tmp;
  wire unequal_tmp;
  wire for_for_for_1_nor_dfs;
  wire [6:0] for_for_row_6_0_lpi_1_dfm;
  wire for_for_for_1_and_2_m1c;
  wire exit_for_for_lpi_1_dfm_5;
  wire for_for_for_1_and_10_m1c;
  wire WX_if_1_and_stg_2_0_sva_mx0;
  wire WX_if_1_and_stg_1_3_sva_mx0;
  wire WX_if_1_and_stg_1_2_sva_mx0;
  wire WX_if_1_and_stg_1_1_sva_mx0;
  wire WX_unequal_tmp_1;
  wire WX_if_1_and_stg_1_0_sva_mx0w0;
  wire for_for_for_1_or_cse;
  wire exit_WY_lpi_1_dfm_2;
  wire [1:0] WX_wx_1_0_lpi_1_dfm;
  wire [2:0] WX_if_1_acc_1_ncse;
  wire [3:0] nl_WX_if_1_acc_1_ncse;
  wire [1:0] WY_wy_1_0_lpi_1_dfm;
  wire for_for_for_1_and_97_cse;
  wire exitL_exit_COL_1_COMP_lpi_1_dfm;
  wire for_for_for_1_asn_rgt_4;
  wire for_for_for_1_for_for_for_1_nor_m1c;
  wire WX_acc_tmp_1;
  wire WY_acc_tmp_1;
  reg reg_output_rsci_oswt_cse;
  reg reg_weight_rsci_oswt_cse;
  reg reg_input_rsci_oswt_cse;
  wire COMP_i_and_cse;
  wire or_79_cse;
  wire WX_if_1_and_cse;
  wire [1:0] WY_mux_3_cse;
  wire nor_41_cse;
  wire or_71_cse;
  wire [1:0] WY_wy_1_0_sva_1;
  wire [2:0] nl_WY_wy_1_0_sva_1;
  wire or_178_tmp;
  wire for_for_for_1_and_285_tmp;
  wire or_tmp_84;
  wire not_tmp_131;
  wire or_tmp_250;
  wire and_119_rgt;
  wire for_for_for_1_and_279_rgt;
  wire [3:0] for_for_for_1_k_mux_itm;
  reg reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_itm;
  reg [2:0] reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_1_itm;
  wire and_235_itm;
  wire [15:0] PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_itm;
  wire [15:0] COL_16_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_15_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_14_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_13_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_12_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_11_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_10_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_9_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_8_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_7_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_6_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_5_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_4_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_3_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_2_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [15:0] COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  wire [1023:0] for_for_out_stencil_value_sva_1_mx0w0;
  wire [1:0] WX_wx_1_0_sva_1;
  wire [2:0] nl_WX_wx_1_0_sva_1;
  wire COMP_i_0_1_lpi_1_dfm;
  wire COMP_i_0_2_lpi_1_dfm;
  wire COMP_i_0_3_lpi_1_dfm;
  wire COMP_i_0_4_lpi_1_dfm;
  wire COMP_i_0_5_lpi_1_dfm;
  wire COMP_i_0_6_lpi_1_dfm;
  wire COMP_i_0_7_lpi_1_dfm;
  wire COMP_i_0_8_lpi_1_dfm;
  wire COMP_i_0_9_lpi_1_dfm;
  wire COMP_i_0_10_lpi_1_dfm;
  wire COMP_i_0_11_lpi_1_dfm;
  wire COMP_i_0_12_lpi_1_dfm;
  wire COMP_i_0_13_lpi_1_dfm;
  wire COMP_i_0_14_lpi_1_dfm;
  wire COMP_i_0_15_lpi_1_dfm;
  wire COMP_i_0_lpi_1_dfm;
  wire exit_for_lpi_1_dfm_3;
  wire [31:0] out_tmp_value_15_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_15_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_14_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_14_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_13_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_13_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_12_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_12_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_11_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_11_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_10_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_10_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_9_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_9_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_8_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_8_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_7_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_7_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_6_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_6_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_5_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_5_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_4_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_4_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_3_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_3_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_2_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_2_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_1_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_1_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_0_31_0_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_0_63_32_lpi_1_mx0w0;
  wire [31:0] out_tmp_value_15_31_0_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_15_63_32_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_14_31_0_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_14_63_32_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_13_31_0_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_13_63_32_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_12_31_0_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_12_63_32_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_11_31_0_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_11_63_32_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_10_31_0_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_10_63_32_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_9_31_0_lpi_1_dfm;
  wire [31:0] out_tmp_value_9_63_32_lpi_1_dfm;
  wire [31:0] out_tmp_value_8_31_0_lpi_1_dfm;
  wire [31:0] out_tmp_value_8_63_32_lpi_1_dfm;
  wire [31:0] out_tmp_value_7_31_0_lpi_1_dfm;
  wire [31:0] out_tmp_value_7_63_32_lpi_1_dfm;
  wire [31:0] out_tmp_value_6_31_0_lpi_1_dfm;
  wire [31:0] out_tmp_value_6_63_32_lpi_1_dfm;
  wire [31:0] out_tmp_value_5_31_0_lpi_1_dfm;
  wire [31:0] out_tmp_value_5_63_32_lpi_1_dfm;
  wire [31:0] out_tmp_value_4_31_0_lpi_1_dfm;
  wire [31:0] out_tmp_value_4_63_32_lpi_1_dfm;
  wire [31:0] out_tmp_value_3_31_0_lpi_1_dfm;
  wire [31:0] out_tmp_value_3_63_32_lpi_1_dfm;
  wire [31:0] out_tmp_value_2_31_0_lpi_1_dfm;
  wire [31:0] out_tmp_value_2_63_32_lpi_1_dfm;
  wire [31:0] out_tmp_value_1_31_0_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_1_63_32_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_0_31_0_lpi_1_dfm_mx0w0;
  wire [31:0] out_tmp_value_0_63_32_lpi_1_dfm_mx0w0;
  wire [31:0] pe_y_reg_value_15_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_15_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_14_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_14_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_13_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_13_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_12_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_12_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_11_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_11_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_10_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_10_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_9_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_9_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_8_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_8_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_7_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_7_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_6_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_6_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_5_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_5_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_4_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_4_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_3_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_3_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_2_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_2_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_1_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_1_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_0_63_32_sva_1_mx0;
  wire [31:0] pe_y_reg_value_0_31_0_sva_1_mx0;
  wire [31:0] pe_y_reg_value_15_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_16_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_16_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_15_31_0_lpi_1_dfm_mx0;
  wire [15:0] in_tmp_16_lpi_1_dfm_1;
  wire [31:0] pe_y_reg_value_14_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_15_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_15_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_14_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_13_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_14_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_14_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_13_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_12_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_13_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_13_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_12_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_11_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_12_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_12_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_11_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_10_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_11_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_11_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_10_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_9_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_10_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_10_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_9_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_8_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_9_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_9_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_8_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_7_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_8_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_8_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_7_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_6_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_7_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_7_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_6_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_5_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_6_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_6_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_5_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_4_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_5_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_5_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_4_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_3_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_4_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_4_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_3_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_2_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_3_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_3_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_2_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_1_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_2_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_2_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_1_31_0_lpi_1_dfm_mx0;
  wire [31:0] pe_y_reg_value_0_63_32_lpi_1_dfm_mx0;
  wire [15:0] COL_1_COMP_tmp_acc_psp_sva;
  wire [16:0] nl_COL_1_COMP_tmp_acc_psp_sva;
  wire [31:0] pe_y_reg_value_0_31_0_lpi_1_dfm_mx0;
  wire [15:0] pe_x_reg_0_lpi_1_dfm;
  wire [1:0] for_ko_2_0_lpi_1_dfm_1_0;
  wire WX_and_16_psp_mx0w0;
  wire WX_and_14_psp_mx0w0;
  wire WX_and_12_psp_mx0w0;
  wire WX_and_10_psp_mx0w0;
  wire WX_and_8_psp_mx0w0;
  wire WX_and_6_psp_mx0w0;
  wire WX_and_4_psp_mx0w0;
  wire WX_and_2_psp_mx0w0;
  wire WX_and_psp_mx0w0;
  wire [15:0] in_tmp_14_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_13_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_12_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_11_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_10_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_9_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_8_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_7_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_6_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_5_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_4_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_3_lpi_1_dfm_1_mx0;
  wire [15:0] in_tmp_2_lpi_1_dfm_1_mx0;
  wire WX_if_1_and_stg_1_1_sva_mx0w0;
  wire WX_if_1_and_stg_1_2_sva_mx0w0;
  wire WX_if_1_and_stg_1_3_sva_mx0w0;
  wire WX_if_1_and_stg_2_0_sva_mx0w0;
  wire [2:0] WX_if_1_acc_decb_sva_3_1_mx0w0;
  wire [3:0] nl_WX_if_1_acc_decb_sva_3_1_mx0w0;
  wire asn_259;
  wire for_for_for_1_asn_426;
  wire for_for_for_1_asn_428;
  wire for_for_for_1_asn_430;
  wire for_for_for_1_asn_432;
  wire asn_261;
  reg reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp;
  reg [2:0] reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp_1;
  wire pe_y_reg_value_and_cse;
  wire PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_and_cse;
  wire for_for_for_1_and_291_cse;
  wire nor_317_cse;
  wire mux_273_cse;
  wire or_395_cse;
  wire and_729_cse;
  wire out_tmp_value_and_26_cse;
  wire for_for_for_1_and_293_cse;
  wire for_for_for_1_and_289_cse;
  wire for_for_row_and_1_cse;
  wire WX_and_19_cse;
  wire for_for_row_and_cse;
  wire for_for_for_1_and_299_cse;
  wire in_tmp_and_1_cse;
  wire pe_x_reg_and_cse;
  wire in_tmp_and_14_cse;
  wire for_for_for_1_and_300_cse;
  wire WY_wy_and_cse;
  wire COL_and_cse;
  wire nand_75_cse;
  wire out_tmp_value_and_1_cse;
  wire out_tmp_value_and_2_cse;
  wire mux_272_cse;
  wire weight_buf_value_and_12_cse;
  wire out_tmp_value_and_25_cse;
  wire weight_buf_value_and_cse;
  wire weight_buf_value_and_2_cse;
  wire weight_buf_value_and_4_cse;
  wire weight_buf_value_and_6_cse;
  wire weight_buf_value_and_8_cse;
  wire weight_buf_value_and_10_cse;
  wire weight_buf_value_and_14_cse;
  wire weight_buf_value_and_16_cse;
  wire [15:0] mux_414_cse;
  wire and_741_tmp;
  wire and_742_tmp;
  wire and_743_tmp;
  wire and_744_tmp;
  wire and_745_tmp;
  wire and_746_tmp;
  wire and_747_tmp;
  wire and_748_tmp;
  wire and_749_tmp;

  wire[0:0] mux_150_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] or_7_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] or_11_nl;
  wire[3:0] WY_WY_and_2_nl;
  wire[0:0] WY_not_10_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] nor_60_nl;
  wire[0:0] nor_61_nl;
  wire[0:0] or_170_nl;
  wire[0:0] WY_WY_and_3_nl;
  wire[0:0] and_55_nl;
  wire[0:0] for_for_for_1_mux1h_196_nl;
  wire[0:0] for_for_for_1_mux1h_193_nl;
  wire[1:0] mux_203_nl;
  wire[0:0] and_241_nl;
  wire[0:0] nor_64_nl;
  wire[0:0] for_for_for_1_nand_nl;
  wire[0:0] for_for_for_1_and_nl;
  wire[0:0] for_for_for_1_and_166_nl;
  wire[31:0] and_59_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] nand_10_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] or_202_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] and_259_nl;
  wire[0:0] nor_315_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] nor_316_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] and_264_nl;
  wire[0:0] nor_312_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] nor_313_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] and_269_nl;
  wire[0:0] nor_309_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] nor_310_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] and_274_nl;
  wire[0:0] nor_306_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] nor_307_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] and_279_nl;
  wire[0:0] nor_303_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] nor_304_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] and_284_nl;
  wire[0:0] nor_300_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] nor_301_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] and_289_nl;
  wire[0:0] nor_297_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] nor_298_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] and_294_nl;
  wire[0:0] nor_294_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] nor_295_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] and_299_nl;
  wire[0:0] nor_291_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] nor_292_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] and_304_nl;
  wire[0:0] nor_288_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] nor_289_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] and_309_nl;
  wire[0:0] nor_285_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] nor_286_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] and_314_nl;
  wire[0:0] nor_282_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] nor_283_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] and_319_nl;
  wire[0:0] nor_279_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] nor_280_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] and_324_nl;
  wire[0:0] nor_276_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] nor_277_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] and_329_nl;
  wire[0:0] nor_273_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] nor_274_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] and_334_nl;
  wire[0:0] nor_270_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] nor_271_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] and_339_nl;
  wire[0:0] nor_267_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] nor_268_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] and_344_nl;
  wire[0:0] nor_264_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] nor_265_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] and_349_nl;
  wire[0:0] nor_261_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] nor_262_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] and_354_nl;
  wire[0:0] nor_258_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] nor_259_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] and_359_nl;
  wire[0:0] nor_255_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] nor_256_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] and_364_nl;
  wire[0:0] nor_252_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] nor_253_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] and_369_nl;
  wire[0:0] nor_249_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] nor_250_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] and_374_nl;
  wire[0:0] nor_246_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] nor_247_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] and_379_nl;
  wire[0:0] nor_243_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] nor_244_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] and_384_nl;
  wire[0:0] nor_240_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] nor_241_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] and_389_nl;
  wire[0:0] nor_237_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] nor_238_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] and_394_nl;
  wire[0:0] nor_234_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] nor_235_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] and_399_nl;
  wire[0:0] nor_231_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] nor_232_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] and_404_nl;
  wire[0:0] nor_228_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] nor_229_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] and_409_nl;
  wire[0:0] nor_225_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] nor_226_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] and_414_nl;
  wire[0:0] nor_222_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] nor_223_nl;
  wire[0:0] and_730_nl;
  wire[0:0] nor_221_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] nor_220_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] and_418_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] nor_217_nl;
  wire[31:0] and_89_nl;
  wire[31:0] and_88_nl;
  wire[31:0] and_87_nl;
  wire[31:0] and_86_nl;
  wire[31:0] and_85_nl;
  wire[31:0] and_84_nl;
  wire[31:0] and_83_nl;
  wire[31:0] and_82_nl;
  wire[31:0] and_81_nl;
  wire[31:0] and_80_nl;
  wire[31:0] and_79_nl;
  wire[31:0] and_78_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] nor_51_nl;
  wire[31:0] and_61_nl;
  wire[31:0] and_60_nl;
  wire[31:0] and_58_nl;
  wire[15:0] mux1h_nl;
  wire[0:0] nor_321_nl;
  wire[0:0] and_751_nl;
  wire[15:0] mux1h_38_nl;
  wire[0:0] nor_322_nl;
  wire[0:0] and_753_nl;
  wire[15:0] mux1h_39_nl;
  wire[0:0] nor_323_nl;
  wire[0:0] and_755_nl;
  wire[15:0] mux1h_40_nl;
  wire[0:0] nor_324_nl;
  wire[0:0] and_757_nl;
  wire[15:0] mux1h_41_nl;
  wire[0:0] nor_325_nl;
  wire[0:0] and_759_nl;
  wire[15:0] mux1h_42_nl;
  wire[0:0] nor_326_nl;
  wire[0:0] and_761_nl;
  wire[15:0] mux1h_43_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] and_763_nl;
  wire[15:0] mux1h_44_nl;
  wire[0:0] nor_328_nl;
  wire[0:0] and_765_nl;
  wire[15:0] mux1h_45_nl;
  wire[0:0] nor_329_nl;
  wire[0:0] and_767_nl;
  wire[0:0] or_68_nl;
  wire[0:0] or_66_nl;
  wire[2:0] WX_if_1_mux_29_nl;
  wire[0:0] and_234_nl;
  wire[0:0] or_75_nl;
  wire[0:0] and_228_nl;
  wire[0:0] and_232_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] nor_39_nl;
  wire[0:0] nor_40_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] nor_35_nl;
  wire[0:0] nor_36_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] nor_31_nl;
  wire[0:0] nor_32_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] nor_27_nl;
  wire[0:0] nor_28_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] nor_23_nl;
  wire[0:0] nor_24_nl;
  wire[0:0] mux_186_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] nor_19_nl;
  wire[0:0] nor_20_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] nor_15_nl;
  wire[0:0] nor_16_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] mux_193_nl;
  wire[0:0] nor_11_nl;
  wire[0:0] nor_12_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] nor_7_nl;
  wire[0:0] nor_8_nl;
  wire[0:0] and_233_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] nor_45_nl;
  wire[0:0] nor_46_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] nor_44_nl;
  wire[0:0] mux_164_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] or_51_nl;
  wire[0:0] or_50_nl;
  wire[0:0] WY_mux_1_nl;
  wire[0:0] nor_63_nl;
  wire[31:0] and_52_nl;
  wire[31:0] and_51_nl;
  wire[31:0] and_50_nl;
  wire[31:0] and_49_nl;
  wire[31:0] and_48_nl;
  wire[31:0] and_47_nl;
  wire[31:0] and_46_nl;
  wire[31:0] and_45_nl;
  wire[31:0] and_44_nl;
  wire[31:0] and_43_nl;
  wire[31:0] and_42_nl;
  wire[31:0] and_41_nl;
  wire[31:0] and_40_nl;
  wire[31:0] and_39_nl;
  wire[31:0] and_38_nl;
  wire[31:0] and_37_nl;
  wire[31:0] and_36_nl;
  wire[31:0] and_35_nl;
  wire[31:0] and_34_nl;
  wire[31:0] and_33_nl;
  wire[31:0] and_32_nl;
  wire[31:0] and_31_nl;
  wire[31:0] and_30_nl;
  wire[31:0] and_29_nl;
  wire[31:0] and_28_nl;
  wire[31:0] and_27_nl;
  wire[31:0] and_26_nl;
  wire[31:0] and_25_nl;
  wire[31:0] and_24_nl;
  wire[31:0] and_23_nl;
  wire[31:0] and_22_nl;
  wire[31:0] and_21_nl;
  wire[31:0] out_tmp_value_mux_nl;
  wire[31:0] out_tmp_value_mux_1_nl;
  wire[31:0] out_tmp_value_mux_2_nl;
  wire[31:0] out_tmp_value_mux_3_nl;
  wire[31:0] out_tmp_value_mux_4_nl;
  wire[31:0] out_tmp_value_mux_5_nl;
  wire[31:0] out_tmp_value_mux_6_nl;
  wire[31:0] out_tmp_value_mux_7_nl;
  wire[31:0] out_tmp_value_mux_8_nl;
  wire[31:0] out_tmp_value_mux_9_nl;
  wire[31:0] out_tmp_value_mux_10_nl;
  wire[31:0] out_tmp_value_mux_11_nl;
  wire[31:0] out_tmp_value_mux_12_nl;
  wire[31:0] out_tmp_value_mux_13_nl;
  wire[31:0] out_tmp_value_mux_14_nl;
  wire[31:0] out_tmp_value_mux_15_nl;
  wire[31:0] out_tmp_value_mux_16_nl;
  wire[31:0] out_tmp_value_mux_17_nl;
  wire[31:0] out_tmp_value_mux_18_nl;
  wire[31:0] out_tmp_value_mux_19_nl;
  wire[31:0] out_tmp_value_mux_20_nl;
  wire[31:0] out_tmp_value_mux_21_nl;
  wire[31:0] out_tmp_value_mux_22_nl;
  wire[31:0] out_tmp_value_mux_23_nl;
  wire[31:0] out_tmp_value_mux_24_nl;
  wire[31:0] out_tmp_value_mux_25_nl;
  wire[31:0] out_tmp_value_mux_26_nl;
  wire[31:0] out_tmp_value_mux_27_nl;
  wire[31:0] out_tmp_value_mux_28_nl;
  wire[31:0] out_tmp_value_mux_29_nl;
  wire[31:0] out_tmp_value_mux_30_nl;
  wire[31:0] out_tmp_value_mux_31_nl;
  wire[15:0] COL_16_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_16_COMP_tmp_mul_nl;
  wire[15:0] COL_15_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_15_COMP_tmp_mul_nl;
  wire[15:0] COL_14_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_14_COMP_tmp_mul_nl;
  wire[15:0] COL_13_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_13_COMP_tmp_mul_nl;
  wire[15:0] COL_12_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_12_COMP_tmp_mul_nl;
  wire[15:0] COL_11_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_11_COMP_tmp_mul_nl;
  wire[15:0] COL_10_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_10_COMP_tmp_mul_nl;
  wire[15:0] COL_9_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_9_COMP_tmp_mul_nl;
  wire[15:0] COL_8_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_8_COMP_tmp_mul_nl;
  wire[15:0] COL_7_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_7_COMP_tmp_mul_nl;
  wire[15:0] COL_6_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_6_COMP_tmp_mul_nl;
  wire[15:0] COL_5_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_5_COMP_tmp_mul_nl;
  wire[15:0] COL_4_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_4_COMP_tmp_mul_nl;
  wire[15:0] COL_3_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_3_COMP_tmp_mul_nl;
  wire[15:0] COL_2_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_2_COMP_tmp_mul_nl;
  wire[15:0] COL_1_COMP_tmp_mul_nl;
  wire signed [32:0] nl_COL_1_COMP_tmp_mul_nl;
  wire[0:0] for_not_39_nl;
  wire[0:0] WX_if_1_mux_26_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] nor_53_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] or_41_nl;
  wire[0:0] or_38_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[31:0] PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_mux_nl;
  wire[31:0] PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_mux_1_nl;
  wire [63:0] nl_PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_rg_a;
  assign PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_mux_nl = MUX_v_32_16_2(pe_y_reg_value_0_63_32_lpi_2,
      pe_y_reg_value_1_63_32_lpi_2, pe_y_reg_value_2_63_32_lpi_2, pe_y_reg_value_3_63_32_lpi_2,
      pe_y_reg_value_4_63_32_lpi_2, pe_y_reg_value_5_63_32_lpi_2, pe_y_reg_value_6_63_32_lpi_2,
      pe_y_reg_value_7_63_32_lpi_2, pe_y_reg_value_8_63_32_lpi_2, pe_y_reg_value_9_63_32_lpi_2,
      pe_y_reg_value_10_63_32_lpi_2, pe_y_reg_value_11_63_32_lpi_2, pe_y_reg_value_12_63_32_lpi_2,
      pe_y_reg_value_13_63_32_lpi_2, pe_y_reg_value_14_63_32_lpi_2, pe_y_reg_value_15_63_32_lpi_2,
      {reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp , reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp_1});
  assign PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_mux_1_nl = MUX_v_32_16_2(pe_y_reg_value_0_31_0_lpi_2,
      pe_y_reg_value_1_31_0_lpi_2, pe_y_reg_value_2_31_0_lpi_2, pe_y_reg_value_3_31_0_lpi_2,
      pe_y_reg_value_4_31_0_lpi_2, pe_y_reg_value_5_31_0_lpi_2, pe_y_reg_value_6_31_0_lpi_2,
      pe_y_reg_value_7_31_0_lpi_2, pe_y_reg_value_8_31_0_lpi_2, pe_y_reg_value_9_31_0_lpi_2,
      pe_y_reg_value_10_31_0_lpi_2, pe_y_reg_value_11_31_0_lpi_2, pe_y_reg_value_12_31_0_lpi_2,
      pe_y_reg_value_13_31_0_lpi_2, pe_y_reg_value_14_31_0_lpi_2, pe_y_reg_value_15_31_0_lpi_2,
      {reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp , reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp_1});
  assign nl_PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_rg_a = {(PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_mux_nl)
      , (PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_mux_1_nl)};
  wire [5:0] nl_PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_rg_s;
  assign nl_PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_rg_s = {PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_lo_conc_1_itm_2_5_1
      , 5'b0};
  wire [63:0] nl_COL_16_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_16_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_15_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_15_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_16_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_16_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_15_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_15_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_14_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_14_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_15_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_15_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_15_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_14_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_14_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_13_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_13_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_14_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_14_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_14_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_13_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_13_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_12_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_12_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_13_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_13_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_13_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_12_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_12_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_11_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_11_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_12_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_12_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_12_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_11_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_11_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_10_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_10_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_11_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_11_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_11_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_10_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_10_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_9_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_9_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_10_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_10_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_10_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_9_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_9_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_8_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_8_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_9_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_9_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_9_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_8_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_8_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_7_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_7_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_8_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_8_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_8_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_7_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_7_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_6_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_6_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_7_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_7_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_7_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_6_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_6_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_5_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_5_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_6_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_6_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_6_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_5_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_5_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_4_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_4_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_5_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_5_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_5_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_4_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_4_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_3_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_3_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_4_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_4_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_4_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_3_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_3_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_2_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_2_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_3_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_3_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_3_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_2_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_2_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_1_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_1_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_2_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_2_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_2_lpi_1_dfm_6
      , 5'b0};
  wire [63:0] nl_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a;
  assign nl_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a = {pe_y_reg_value_0_63_32_lpi_1_dfm_mx0
      , pe_y_reg_value_0_31_0_lpi_1_dfm_mx0};
  wire [5:0] nl_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s;
  assign nl_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s = {COMP_i_0_1_lpi_1_dfm_6
      , 5'b0};
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_rg (
      .a(nl_PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_rg_a[63:0]),
      .s(nl_PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_rg_s[5:0]),
      .z(PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_16_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg
      (
      .a(nl_COL_16_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_16_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_16_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_15_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg
      (
      .a(nl_COL_15_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_15_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_15_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_14_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg
      (
      .a(nl_COL_14_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_14_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_14_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_13_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg
      (
      .a(nl_COL_13_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_13_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_13_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_12_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg
      (
      .a(nl_COL_12_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_12_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_12_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_11_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg
      (
      .a(nl_COL_11_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_11_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_11_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_10_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg
      (
      .a(nl_COL_10_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_10_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_10_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_9_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg (
      .a(nl_COL_9_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_9_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_9_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_8_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg (
      .a(nl_COL_8_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_8_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_8_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_7_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg (
      .a(nl_COL_7_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_7_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_7_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_6_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg (
      .a(nl_COL_6_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_6_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_6_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_5_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg (
      .a(nl_COL_5_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_5_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_5_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_4_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg (
      .a(nl_COL_4_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_4_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_4_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_3_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg (
      .a(nl_COL_3_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_3_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_3_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_2_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg (
      .a(nl_COL_2_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_2_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_2_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  mgc_shift_r_v4 #(.width_a(32'sd64),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd16)) COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg (
      .a(nl_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_a[63:0]),
      .s(nl_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_rg_s[5:0]),
      .z(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm)
    );
  systolic_array_core_input_rsci systolic_array_core_input_rsci_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_z(input_rsc_z),
      .input_rsc_vz(input_rsc_vz),
      .input_rsc_lz(input_rsc_lz),
      .core_wen(core_wen),
      .input_rsci_oswt(reg_input_rsci_oswt_cse),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .input_rsci_d_mxwt(input_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  systolic_array_core_weight_rsci systolic_array_core_weight_rsci_inst (
      .clk(clk),
      .rst(rst),
      .weight_rsc_z(weight_rsc_z),
      .weight_rsc_vz(weight_rsc_vz),
      .weight_rsc_lz(weight_rsc_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .weight_rsci_oswt(reg_weight_rsci_oswt_cse),
      .weight_rsci_wen_comp(weight_rsci_wen_comp),
      .weight_rsci_d_mxwt(weight_rsci_d_mxwt)
    );
  systolic_array_core_output_rsci systolic_array_core_output_rsci_inst (
      .clk(clk),
      .rst(rst),
      .output_rsc_z(output_rsc_z),
      .output_rsc_vz(output_rsc_vz),
      .output_rsc_lz(output_rsc_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .output_rsci_oswt(reg_output_rsci_oswt_cse),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .output_rsci_d(output_rsci_d)
    );
  systolic_array_core_staller systolic_array_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .core_wten(core_wten),
      .weight_rsci_wen_comp(weight_rsci_wen_comp),
      .output_rsci_wen_comp(output_rsci_wen_comp)
    );
  assign for_for_for_1_and_289_cse = core_wen & main_stage_0_2 & (~ lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign or_7_nl = (~((~ exit_for_for_for_1_lpi_1_dfm_1_st_3) | lfst_exit_for_for_for_1_lpi_1_dfm_st_1_0))
      | for_for_for_1_equal_tmp_2;
  assign mux_148_nl = MUX_s_1_2_2(mux_tmp, or_tmp_5, or_7_nl);
  assign or_11_nl = (~ exitL_exit_COL_1_COMP_lpi_1_dfm_4) | for_for_for_1_equal_tmp_2;
  assign mux_149_nl = MUX_s_1_2_2(mux_tmp, or_tmp_5, or_11_nl);
  assign mux_150_nl = MUX_s_1_2_2((mux_149_nl), (mux_148_nl), lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign pe_y_reg_value_and_cse = core_wen & (~((~ main_stage_0_3) | for_for_for_1_equal_tmp_10
      | for_for_for_1_equal_tmp_12)) & (mux_150_nl);
  assign PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_and_cse = core_wen & (for_for_for_1_equal_tmp_2
      | exit_for_for_for_1_lpi_1_dfm_1_st_3) & main_stage_0_2 & and_dcpl_1;
  assign for_for_for_1_and_291_cse = core_wen & main_stage_0_2;
  assign for_for_row_and_cse = core_wen & or_tmp_4;
  assign COMP_i_and_cse = core_wen & (~ and_dcpl_65);
  assign WY_wy_and_cse = core_wen & for_for_for_1_nand_2_tmp;
  assign for_for_row_and_1_cse = core_wen & or_dcpl_15;
  assign nor_317_cse = ~((~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4)
      | for_for_for_1_nor_dfs_7 | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign and_730_nl = lfst_exit_for_for_1_lpi_1_dfm_1 & main_stage_0_4;
  assign nor_221_nl = ~((~ lfst_exit_for_for_1_lpi_2) | exitL_exit_for_sva | exit_for_lpi_1_dfm_4
      | (~ main_stage_0_4));
  assign mux_273_cse = MUX_s_1_2_2((nor_221_nl), (and_730_nl), main_stage_0_2);
  assign or_395_cse = (~ main_stage_0_2) | lfst_exit_for_for_1_lpi_1_dfm_1;
  assign and_729_cse = lfst_exit_for_for_for_1_lpi_1_dfm_9_1_1 & for_for_for_1_equal_tmp_10;
  assign nor_220_nl = ~((~ unequal_tmp_6) | COMP_and_13_mdf_sva_6 | (~(for_for_for_1_nor_dfs_6
      & or_tmp_250)));
  assign mux_271_nl = MUX_s_1_2_2((nor_220_nl), or_tmp_250, and_729_cse);
  assign mux_272_cse = MUX_s_1_2_2((mux_271_nl), or_tmp_250, for_for_for_1_equal_tmp_12);
  assign and_418_nl = or_395_cse & mux_272_cse;
  assign mux_274_nl = MUX_s_1_2_2(mux_273_cse, (and_418_nl), main_stage_0_3);
  assign out_tmp_value_and_1_cse = (mux_274_nl) & core_wen;
  assign nand_75_cse = ~(for_for_for_1_equal_tmp_10 & ((~ for_for_row_6_0_lpi_1_dfm_6_6_1)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | for_for_for_1_nor_dfs_7 | for_for_for_1_equal_tmp_11
      | for_for_for_1_equal_tmp_13 | (~ main_stage_0_4)));
  assign nor_217_nl = ~((~((~ main_stage_0_2) | lfst_exit_for_for_1_lpi_1_dfm_1))
      | lfst_exit_for_for_for_1_lpi_1_dfm_9_1_1 | nand_75_cse);
  assign mux_276_nl = MUX_s_1_2_2(mux_273_cse, (nor_217_nl), main_stage_0_3);
  assign out_tmp_value_and_2_cse = (mux_276_nl) & core_wen;
  assign nor_51_nl = ~((~ unequal_tmp_6) | COMP_and_13_mdf_sva_6 | (~(for_for_for_1_nor_dfs_6
      & or_395_cse)));
  assign mux_154_nl = MUX_s_1_2_2((nor_51_nl), or_395_cse, and_729_cse);
  assign mux_155_nl = MUX_s_1_2_2((mux_154_nl), or_395_cse, for_for_for_1_equal_tmp_12);
  assign out_tmp_value_and_25_cse = mux_272_cse & main_stage_0_3 & core_wen & (mux_155_nl);
  assign out_tmp_value_and_26_cse = (for_for_for_1_equal_tmp_13 | for_for_for_1_equal_tmp_11
      | for_for_for_1_nor_dfs_7 | (~(main_stage_0_4 & lfst_exit_for_for_1_lpi_1_dfm_4
      & for_for_row_6_0_lpi_1_dfm_6_6_1))) & for_for_for_1_equal_tmp_10 & core_wen
      & or_395_cse & (~ lfst_exit_for_for_for_1_lpi_1_dfm_9_1_1) & main_stage_0_3;
  assign for_for_for_1_and_293_cse = core_wen & or_395_cse & main_stage_0_3;
  assign and_741_tmp = WX_and_16_psp_mx0w0 & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign and_742_tmp = WX_and_14_psp_mx0w0 & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign and_743_tmp = WX_and_12_psp_mx0w0 & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign and_744_tmp = WX_and_10_psp_mx0w0 & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign and_745_tmp = WX_and_8_psp_mx0w0 & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign and_746_tmp = WX_and_6_psp_mx0w0 & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign and_747_tmp = WX_and_4_psp_mx0w0 & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign and_748_tmp = WX_and_2_psp_mx0w0 & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign and_749_tmp = WX_and_psp_mx0w0 & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign or_66_nl = or_dcpl_38 | WY_acc_tmp_1;
  assign WY_mux_3_cse = MUX_v_2_2_2(2'b10, 2'b1, or_66_nl);
  assign for_for_for_1_and_299_cse = core_wen & or_71_cse;
  assign or_71_cse = or_dcpl_7 | (~ lfst_exit_for_for_1_lpi_2) | (~ lfst_exit_for_for_for_1_lpi_1_1_1);
  assign and_234_nl = lfst_exit_for_for_1_lpi_1_dfm & and_dcpl_59;
  assign WX_if_1_mux_29_nl = MUX_v_3_2_2(WX_if_1_acc_decb_sva_3_1_mx0w0, pref_pref_pref_6_3_0_1_lpi_1_3_1_1,
      and_234_nl);
  assign for_for_for_1_k_mux_itm = MUX_v_4_2_2(for_for_for_1_k_4_0_lpi_1_3_0_1, ({1'b0
      , (WX_if_1_mux_29_nl)}), or_71_cse);
  assign nor_41_cse = ~((~((~ lfst_exit_for_for_for_1_lpi_1_0_1) | exitL_exit_COL_1_COMP_lpi_1
      | (~ lfst_exit_WX_1_lpi_1))) | lfst_exit_for_for_for_1_lpi_1_1_1);
  assign or_79_cse = (for_for_row_slc_for_for_row_6_0_5_0_1_itm_3!=6'b000000);
  assign nor_39_nl = ~((~ WX_if_1_and_stg_1_1_sva) | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b01)
      | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign nor_40_nl = ~((WX_if_1_acc_decb_sva_1_3_1_1[0]) | (~ out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1)
      | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b01) | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign mux_165_nl = MUX_s_1_2_2((nor_40_nl), (nor_39_nl), or_79_cse);
  assign mux_166_nl = MUX_s_1_2_2((mux_165_nl), WX_and_11_psp_1, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign weight_buf_value_and_cse = core_wen & (~((~ (mux_166_nl)) | or_dcpl_51));
  assign nor_35_nl = ~((~ WX_if_1_and_stg_1_1_sva) | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b00)
      | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign nor_36_nl = ~((WX_if_1_acc_decb_sva_1_3_1_1[0]) | (~ out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1)
      | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b00) | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign mux_169_nl = MUX_s_1_2_2((nor_36_nl), (nor_35_nl), or_79_cse);
  assign mux_170_nl = MUX_s_1_2_2((mux_169_nl), WX_and_3_psp_1, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign weight_buf_value_and_2_cse = core_wen & (~((~ (mux_170_nl)) | or_dcpl_51));
  assign nor_31_nl = ~((~ WX_if_1_and_stg_1_2_sva) | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b01)
      | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign nor_32_nl = ~((~ (WX_if_1_acc_decb_sva_1_3_1_1[0])) | out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1
      | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b01) | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign mux_173_nl = MUX_s_1_2_2((nor_32_nl), (nor_31_nl), or_79_cse);
  assign mux_174_nl = MUX_s_1_2_2((mux_173_nl), WX_and_13_psp_1, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign weight_buf_value_and_4_cse = core_wen & (~((~ (mux_174_nl)) | or_dcpl_51));
  assign nor_27_nl = ~((~ WX_if_1_and_stg_1_2_sva) | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b00)
      | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign nor_28_nl = ~((~ (WX_if_1_acc_decb_sva_1_3_1_1[0])) | out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1
      | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b00) | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign mux_177_nl = MUX_s_1_2_2((nor_28_nl), (nor_27_nl), or_79_cse);
  assign mux_178_nl = MUX_s_1_2_2((mux_177_nl), WX_and_5_psp_1, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign weight_buf_value_and_6_cse = core_wen & (~((~ (mux_178_nl)) | or_dcpl_51));
  assign nor_23_nl = ~((~ WX_if_1_and_stg_1_3_sva) | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b01)
      | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign nor_24_nl = ~((~ (WX_if_1_acc_decb_sva_1_3_1_1[0])) | (~ out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1)
      | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b01) | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign mux_181_nl = MUX_s_1_2_2((nor_24_nl), (nor_23_nl), or_79_cse);
  assign mux_182_nl = MUX_s_1_2_2((mux_181_nl), WX_and_15_psp_1, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign weight_buf_value_and_8_cse = core_wen & (~((~ (mux_182_nl)) | or_dcpl_51));
  assign nor_19_nl = ~((~ WX_if_1_and_stg_1_3_sva) | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b00)
      | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign nor_20_nl = ~((~ (WX_if_1_acc_decb_sva_1_3_1_1[0])) | (~ out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1)
      | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b00) | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign mux_185_nl = MUX_s_1_2_2((nor_20_nl), (nor_19_nl), or_79_cse);
  assign mux_186_nl = MUX_s_1_2_2((mux_185_nl), WX_and_7_psp_1, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign weight_buf_value_and_10_cse = core_wen & (~((~ (mux_186_nl)) | or_dcpl_51));
  assign nor_15_nl = ~((~ WX_if_1_and_stg_2_0_sva) | (~ (WX_if_1_acc_decb_sva_1_3_1_1[2]))
      | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign nor_16_nl = ~((WX_if_1_acc_decb_sva_1_3_1_1[1:0]!=2'b00) | out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1
      | (~ (WX_if_1_acc_decb_sva_1_3_1_1[2])) | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign mux_189_nl = MUX_s_1_2_2((nor_16_nl), (nor_15_nl), or_79_cse);
  assign mux_190_nl = MUX_s_1_2_2((mux_189_nl), WX_and_17_psp_1, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign weight_buf_value_and_12_cse = core_wen & (~((~ (mux_190_nl)) | or_dcpl_51));
  assign nor_11_nl = ~((~ WX_if_1_and_stg_2_0_sva) | (WX_if_1_acc_decb_sva_1_3_1_1[2])
      | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign nor_12_nl = ~((WX_if_1_acc_decb_sva_1_3_1_1[1:0]!=2'b00) | out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1
      | (WX_if_1_acc_decb_sva_1_3_1_1[2]) | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign mux_193_nl = MUX_s_1_2_2((nor_12_nl), (nor_11_nl), or_79_cse);
  assign mux_194_nl = MUX_s_1_2_2((mux_193_nl), WX_and_1_psp_1, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign weight_buf_value_and_14_cse = core_wen & (~((~ (mux_194_nl)) | or_dcpl_51));
  assign nor_7_nl = ~((~ WX_if_1_and_stg_1_0_sva) | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b01)
      | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign nor_8_nl = ~((WX_if_1_acc_decb_sva_1_3_1_1[0]) | out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1
      | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b01) | (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000));
  assign mux_197_nl = MUX_s_1_2_2((nor_8_nl), (nor_7_nl), or_79_cse);
  assign mux_198_nl = MUX_s_1_2_2((mux_197_nl), WX_and_9_psp_1, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign weight_buf_value_and_16_cse = core_wen & (~((~ (mux_198_nl)) | or_dcpl_51));
  assign WX_and_19_cse = core_wen & (~(or_dcpl_70 | lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1))
      & (~ or_tmp_4);
  assign WX_if_1_and_cse = core_wen & (~(or_dcpl_70 | (for_for_row_slc_for_for_row_6_0_5_0_1_itm_3[3])
      | (for_for_row_slc_for_for_row_6_0_5_0_1_itm_3[5]) | (for_for_row_slc_for_for_row_6_0_5_0_1_itm_3[2])
      | or_dcpl_72 | (for_for_row_slc_for_for_row_6_0_5_0_1_itm_3[4]) | lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1));
  assign and_119_rgt = WX_unequal_tmp_5 & exitL_exit_COL_1_COMP_lpi_1_dfm_4 & (~
      for_for_for_1_or_cse) & main_stage_0_2;
  assign in_tmp_and_1_cse = core_wen & (~ or_dcpl_51) & and_dcpl_38;
  assign for_for_for_1_and_279_rgt = COMP_and_13_mdf_sva_5 & (~ for_for_for_1_or_cse)
      & main_stage_0_2;
  assign pe_x_reg_and_cse = core_wen & (~ or_dcpl_51) & and_dcpl_48;
  assign in_tmp_and_14_cse = core_wen & (~(or_dcpl_50 | for_for_for_1_equal_tmp_2))
      & and_dcpl_48;
  assign for_for_for_1_and_300_cse = core_wen & lfst_exit_for_lpi_1_dfm & lfst_exit_for_for_1_lpi_2
      & main_stage_0_2;
  assign and_235_itm = lfst_exit_for_for_for_1_lpi_1_1_1 & lfst_exit_for_for_1_lpi_2;
  assign mux_161_nl = MUX_s_1_2_2(and_dcpl_27, or_dcpl_18, COMP_and_13_tmp);
  assign mux_162_nl = MUX_s_1_2_2((~ (mux_161_nl)), or_dcpl_14, WY_mux_6_tmp[1]);
  assign or_51_nl = (~(lfst_exit_for_for_for_1_lpi_1_0_1 | (~ lfst_exit_for_for_for_1_lpi_1_1_1)
      | (~ lfst_exit_for_for_1_lpi_2))) | exitL_exit_for_sva | exit_for_lpi_1_dfm_4;
  assign or_50_nl = (~ (for_for_row_6_0_lpi_3[6])) | (WY_mux_6_tmp[1]);
  assign mux_163_nl = MUX_s_1_2_2((or_51_nl), or_dcpl_18, or_50_nl);
  assign mux_164_nl = MUX_s_1_2_2((~ (mux_163_nl)), (mux_162_nl), WY_mux_6_tmp[0]);
  assign COL_and_cse = core_wen & (~ and_dcpl_63) & (mux_164_nl);
  assign for_for_out_stencil_value_sva_1_mx0w0 = writeslice_1024_5_32(for_for_for_1_asn_itm_2,
      {{16{PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_itm[15]}}, PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_rshift_itm},
      {reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp , reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp_1
      , PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_lo_conc_1_itm_2_5_1}, 32, 0);
  assign lfst_exit_for_for_for_1_lpi_1_dfm_1 = lfst_exit_for_for_for_1_lpi_1_1_1
      & lfst_exit_for_for_1_lpi_1_dfm;
  assign lfst_exit_for_for_for_1_lpi_1_dfm_0 = lfst_exit_for_for_for_1_lpi_1_0_1
      & lfst_exit_for_for_1_lpi_1_dfm;
  assign for_for_row_6_0_lpi_1_dfm = MUX_v_7_2_2(7'b0000000, for_for_row_6_0_lpi_3,
      lfst_exit_for_lpi_1_dfm);
  assign WY_acc_tmp_1 = (WY_wy_1_0_sva_1[0]) ^ (WY_wy_1_0_sva_1[1]);
  assign nl_WY_wy_1_0_sva_1 = WY_wy_1_0_lpi_1_dfm + 2'b1;
  assign WY_wy_1_0_sva_1 = nl_WY_wy_1_0_sva_1[1:0];
  assign WY_wy_1_0_lpi_1_dfm = MUX_v_2_2_2(2'b00, WY_wy_1_0_lpi_3, lfst_exit_for_for_1_lpi_1_dfm);
  assign WX_acc_tmp_1 = (WX_wx_1_0_sva_1[0]) ^ (WX_wx_1_0_sva_1[1]);
  assign nl_WX_wx_1_0_sva_1 = WX_wx_1_0_lpi_1_dfm + 2'b1;
  assign WX_wx_1_0_sva_1 = nl_WX_wx_1_0_sva_1[1:0];
  assign WX_wx_1_0_lpi_1_dfm = MUX_v_2_2_2(2'b00, WX_wx_1_0_lpi_3, WY_unequal_tmp);
  assign WY_mux_1_nl = MUX_s_1_2_2((~ WY_acc_tmp_1), exit_WY_sva_2, or_dcpl_38);
  assign exit_WY_lpi_1_dfm_2 = (WY_mux_1_nl) & exit_WX_lpi_1_dfm_1;
  assign exit_WX_lpi_1_dfm_1 = (~ WX_acc_tmp_1) & COMP_and_13_tmp;
  assign COMP_and_13_tmp = COMP_i_0_1_lpi_1_dfm & COMP_i_0_2_lpi_1_dfm & COMP_i_0_3_lpi_1_dfm
      & COMP_i_0_4_lpi_1_dfm & COMP_i_0_5_lpi_1_dfm & COMP_i_0_6_lpi_1_dfm & COMP_i_0_7_lpi_1_dfm
      & COMP_i_0_8_lpi_1_dfm & COMP_i_0_9_lpi_1_dfm & COMP_i_0_10_lpi_1_dfm & COMP_i_0_11_lpi_1_dfm
      & COMP_i_0_12_lpi_1_dfm & COMP_i_0_13_lpi_1_dfm & COMP_i_0_14_lpi_1_dfm & COMP_i_0_15_lpi_1_dfm
      & COMP_i_0_lpi_1_dfm;
  assign COMP_i_0_1_lpi_1_dfm = COMP_i_0_1_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_2_lpi_1_dfm = COMP_i_0_2_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_3_lpi_1_dfm = COMP_i_0_3_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_4_lpi_1_dfm = COMP_i_0_4_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_5_lpi_1_dfm = COMP_i_0_5_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_6_lpi_1_dfm = COMP_i_0_6_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_7_lpi_1_dfm = COMP_i_0_7_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_8_lpi_1_dfm = COMP_i_0_8_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_9_lpi_1_dfm = COMP_i_0_9_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_10_lpi_1_dfm = COMP_i_0_10_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_11_lpi_1_dfm = COMP_i_0_11_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_12_lpi_1_dfm = COMP_i_0_12_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_13_lpi_1_dfm = COMP_i_0_13_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_14_lpi_1_dfm = COMP_i_0_14_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_15_lpi_1_dfm = COMP_i_0_15_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign COMP_i_0_lpi_1_dfm = COMP_i_0_lpi_1 & (~ exitL_exit_COL_1_COMP_lpi_1_dfm);
  assign exitL_exit_COL_1_COMP_lpi_1_dfm = exitL_exit_COL_1_COMP_lpi_1 | (~(lfst_exit_WX_1_lpi_1
      & WY_unequal_tmp));
  assign WY_unequal_tmp = lfst_exit_for_for_for_1_lpi_1_dfm_1 | lfst_exit_for_for_for_1_lpi_1_dfm_0;
  assign for_for_for_1_for_for_for_1_nor_m1c = ~(exit_WX_lpi_1_dfm_1 | lfst_exit_for_for_for_1_lpi_1_dfm_1);
  assign or_178_tmp = (exit_WX_lpi_1_dfm_1 & (~ lfst_exit_for_for_for_1_lpi_1_dfm_1)
      & (~ WY_acc_tmp_1)) | (COMP_and_13_tmp & for_for_for_1_for_for_for_1_nor_m1c);
  assign for_for_for_1_and_285_tmp = (~ COMP_and_13_tmp) & for_for_for_1_for_for_for_1_nor_m1c;
  assign nor_63_nl = ~(for_for_for_1_and_285_tmp | or_178_tmp);
  assign for_for_for_1_for_for_for_1_for_for_for_1_mux1h_1_tmp = MUX1HOT_v_2_3_2((signext_2_1(~
      WY_acc_tmp_1)), WX_wx_1_0_lpi_1_dfm, WX_wx_1_0_sva_1, {(nor_63_nl) , for_for_for_1_and_285_tmp
      , or_178_tmp});
  assign nl_for_for_acc_1_tmp = conv_u2u_6_7(for_for_row_6_0_lpi_1_dfm[5:0]) + 7'b1;
  assign for_for_acc_1_tmp = nl_for_for_acc_1_tmp[6:0];
  assign nl_for_for_for_1_acc_1_tmp = conv_u2u_4_5(for_for_for_1_k_4_0_lpi_1_3_0_1)
      + 5'b1;
  assign for_for_for_1_acc_1_tmp = nl_for_for_for_1_acc_1_tmp[4:0];
  assign exit_for_for_lpi_1_dfm_5 = (for_for_acc_1_tmp[6]) & exit_for_for_for_1_lpi_1_dfm_1;
  assign exit_for_for_for_1_lpi_1_dfm_1 = (for_for_for_1_acc_1_tmp[4]) & for_for_for_1_for_q_0_lpi_2;
  assign for_for_for_1_asn_rgt_4 = (~ for_for_for_1_for_q_0_lpi_2) & for_for_for_1_equal_tmp;
  assign lfst_exit_for_for_1_lpi_1_dfm = lfst_exit_for_for_1_lpi_2 & lfst_exit_for_lpi_1_dfm;
  assign for_for_for_1_nand_2_tmp = ~(exit_for_for_lpi_1_dfm_5 & for_for_for_1_equal_tmp);
  assign lfst_exit_for_lpi_1_dfm = ~(exit_for_lpi_1_dfm_4 | exitL_exit_for_sva);
  assign exit_for_lpi_1_dfm_3 = (for_acc_2_tmp[2]) & exit_for_for_lpi_1_dfm_5 & for_for_for_1_equal_tmp;
  assign and_52_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_33_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_15_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_52_nl), out_tmp_value_15_31_0_lpi_1_dfm_11,
      COMP_mux_23_itm_2, out_tmp_value_15_31_0_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_51_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_32_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_15_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_51_nl), out_tmp_value_15_63_32_lpi_1_dfm_11,
      COMP_mux_24_itm_2, out_tmp_value_15_63_32_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_50_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_31_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_14_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_50_nl), out_tmp_value_14_31_0_lpi_1_dfm_11,
      COMP_mux_21_itm_2, out_tmp_value_14_31_0_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_49_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_30_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_14_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_49_nl), out_tmp_value_14_63_32_lpi_1_dfm_11,
      COMP_mux_22_itm_2, out_tmp_value_14_63_32_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_48_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_29_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_13_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_48_nl), out_tmp_value_13_31_0_lpi_1_dfm_11,
      COMP_mux_2_itm_2, out_tmp_value_13_31_0_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_47_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_28_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_13_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_47_nl), out_tmp_value_13_63_32_lpi_1_dfm_11,
      COMP_mux_20_itm_2, out_tmp_value_13_63_32_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_46_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_27_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_12_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_46_nl), out_tmp_value_12_31_0_lpi_1_dfm_11,
      COMP_mux_18_itm_2, out_tmp_value_12_31_0_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_45_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_26_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_12_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_45_nl), out_tmp_value_12_63_32_lpi_1_dfm_11,
      COMP_mux_19_itm_2, out_tmp_value_12_63_32_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_44_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_25_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_11_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_44_nl), out_tmp_value_11_31_0_lpi_1_dfm_11,
      COMP_mux_16_itm_2, out_tmp_value_11_31_0_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_43_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_24_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_11_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_43_nl), out_tmp_value_11_63_32_lpi_1_dfm_11,
      COMP_mux_17_itm_2, out_tmp_value_11_63_32_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_42_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_23_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_10_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_42_nl), out_tmp_value_10_31_0_lpi_1_dfm_11,
      COMP_mux_14_itm_2, out_tmp_value_10_31_0_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_41_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_22_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_10_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_41_nl), out_tmp_value_10_63_32_lpi_1_dfm_11,
      COMP_mux_15_itm_2, out_tmp_value_10_63_32_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_40_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_21_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_9_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_40_nl), out_tmp_value_9_31_0_lpi_1_dfm_13,
      COMP_mux_8_itm_2, out_tmp_value_9_31_0_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_39_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_20_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_9_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_39_nl), out_tmp_value_9_63_32_lpi_1_dfm_13,
      COMP_mux_9_itm_2, out_tmp_value_9_63_32_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_38_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_19_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_8_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_38_nl), out_tmp_value_8_31_0_lpi_1_dfm_13,
      COMP_mux_6_itm_2, out_tmp_value_8_31_0_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_37_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_18_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_8_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_37_nl), out_tmp_value_8_63_32_lpi_1_dfm_13,
      COMP_mux_7_itm_2, out_tmp_value_8_63_32_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_36_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_17_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_7_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_36_nl), out_tmp_value_7_31_0_lpi_1_dfm_13,
      COMP_mux_4_itm_2, out_tmp_value_7_31_0_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_35_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_16_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_7_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_35_nl), out_tmp_value_7_63_32_lpi_1_dfm_13,
      COMP_mux_5_itm_2, out_tmp_value_7_63_32_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_34_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_15_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_6_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_34_nl), out_tmp_value_6_31_0_lpi_1_dfm_13,
      COMP_mux_32_itm_2, out_tmp_value_6_31_0_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_33_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_14_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_6_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_33_nl), out_tmp_value_6_63_32_lpi_1_dfm_13,
      COMP_mux_33_itm_2, out_tmp_value_6_63_32_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_32_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_13_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_5_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_32_nl), out_tmp_value_5_31_0_lpi_1_dfm_13,
      COMP_mux_30_itm_2, out_tmp_value_5_31_0_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_31_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_12_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_5_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_31_nl), out_tmp_value_5_63_32_lpi_1_dfm_13,
      COMP_mux_31_itm_2, out_tmp_value_5_63_32_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_30_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_11_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_4_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_30_nl), out_tmp_value_4_31_0_lpi_1_dfm_13,
      COMP_mux_29_itm_2, out_tmp_value_4_31_0_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_29_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_10_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_4_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_29_nl), out_tmp_value_4_63_32_lpi_1_dfm_13,
      COMP_mux_3_itm_2, out_tmp_value_4_63_32_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_28_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_9_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_3_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_28_nl), out_tmp_value_3_31_0_lpi_1_dfm_13,
      COMP_mux_27_itm_2, out_tmp_value_3_31_0_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_27_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_8_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_3_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_27_nl), out_tmp_value_3_63_32_lpi_1_dfm_13,
      COMP_mux_28_itm_2, out_tmp_value_3_63_32_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_26_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_7_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_2_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_26_nl), out_tmp_value_2_31_0_lpi_1_dfm_13,
      COMP_mux_25_itm_2, out_tmp_value_2_31_0_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_25_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_6_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_2_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_25_nl), out_tmp_value_2_63_32_lpi_1_dfm_13,
      COMP_mux_26_itm_2, out_tmp_value_2_63_32_lpi_1_dfm_12, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_24_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_5_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_1_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_24_nl), out_tmp_value_1_31_0_lpi_1_dfm_11,
      COMP_mux_12_itm_2, out_tmp_value_1_31_0_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_23_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_4_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_1_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_23_nl), out_tmp_value_1_63_32_lpi_1_dfm_11,
      COMP_mux_13_itm_2, out_tmp_value_1_63_32_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_22_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_3_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_0_31_0_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_22_nl), out_tmp_value_0_31_0_lpi_1_dfm_10,
      COMP_mux_10_itm_2, out_tmp_value_0_31_0_lpi_2, {for_for_for_1_asn_426 , for_for_for_1_asn_428
      , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign and_21_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, COMP_mux_2_itm_2,
      for_for_row_6_0_lpi_1_dfm_7_6_1);
  assign out_tmp_value_0_63_32_lpi_1_mx0w0 = MUX1HOT_v_32_4_2((and_21_nl), out_tmp_value_0_63_32_lpi_1_dfm_11,
      COMP_mux_11_itm_2, out_tmp_value_0_63_32_lpi_1_dfm_10, {for_for_for_1_asn_426
      , for_for_for_1_asn_428 , for_for_for_1_asn_430 , for_for_for_1_asn_432});
  assign out_tmp_value_mux_nl = MUX_v_32_2_2(out_tmp_value_11_63_32_lpi_1_dfm_10,
      out_tmp_value_15_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_15_31_0_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_1_nl = MUX_v_32_2_2(out_tmp_value_11_63_32_lpi_1_dfm_11,
      out_tmp_value_15_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_15_63_32_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_1_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_2_nl = MUX_v_32_2_2(out_tmp_value_11_31_0_lpi_1_dfm_10,
      out_tmp_value_14_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_14_31_0_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_2_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_3_nl = MUX_v_32_2_2(out_tmp_value_11_31_0_lpi_1_dfm_11,
      out_tmp_value_14_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_14_63_32_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_3_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_4_nl = MUX_v_32_2_2(out_tmp_value_10_63_32_lpi_1_dfm_10,
      out_tmp_value_13_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_13_31_0_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_4_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_5_nl = MUX_v_32_2_2(out_tmp_value_10_63_32_lpi_1_dfm_11,
      out_tmp_value_13_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_13_63_32_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_5_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_6_nl = MUX_v_32_2_2(out_tmp_value_10_31_0_lpi_1_dfm_10,
      out_tmp_value_12_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_12_31_0_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_6_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_7_nl = MUX_v_32_2_2(out_tmp_value_10_31_0_lpi_1_dfm_11,
      out_tmp_value_12_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_12_63_32_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_7_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_8_nl = MUX_v_32_2_2(out_tmp_value_1_63_32_lpi_1_dfm_10,
      out_tmp_value_11_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_11_31_0_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_8_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_9_nl = MUX_v_32_2_2(out_tmp_value_1_63_32_lpi_1_dfm_11,
      out_tmp_value_11_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_11_63_32_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_9_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_10_nl = MUX_v_32_2_2(out_tmp_value_1_31_0_lpi_1_dfm_10,
      out_tmp_value_10_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_10_31_0_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_10_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_11_nl = MUX_v_32_2_2(out_tmp_value_1_31_0_lpi_1_dfm_11,
      out_tmp_value_10_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_10_63_32_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_11_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_12_nl = MUX_v_32_2_2(out_tmp_value_15_63_32_lpi_1_dfm_10,
      out_tmp_value_9_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_9_31_0_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_12_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_13_nl = MUX_v_32_2_2(out_tmp_value_15_63_32_lpi_1_dfm_11,
      out_tmp_value_9_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_9_63_32_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_13_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_14_nl = MUX_v_32_2_2(out_tmp_value_15_31_0_lpi_1_dfm_10,
      out_tmp_value_8_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_8_31_0_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_14_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_15_nl = MUX_v_32_2_2(out_tmp_value_15_31_0_lpi_1_dfm_11,
      out_tmp_value_8_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_8_63_32_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_15_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_16_nl = MUX_v_32_2_2(out_tmp_value_14_63_32_lpi_1_dfm_10,
      out_tmp_value_7_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_7_31_0_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_16_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_17_nl = MUX_v_32_2_2(out_tmp_value_14_63_32_lpi_1_dfm_11,
      out_tmp_value_7_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_7_63_32_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_17_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_18_nl = MUX_v_32_2_2(out_tmp_value_14_31_0_lpi_1_dfm_10,
      out_tmp_value_6_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_6_31_0_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_18_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_19_nl = MUX_v_32_2_2(out_tmp_value_14_31_0_lpi_1_dfm_11,
      out_tmp_value_6_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_6_63_32_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_19_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_20_nl = MUX_v_32_2_2(out_tmp_value_13_63_32_lpi_1_dfm_10,
      out_tmp_value_5_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_5_31_0_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_20_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_21_nl = MUX_v_32_2_2(out_tmp_value_13_63_32_lpi_1_dfm_11,
      out_tmp_value_5_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_5_63_32_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_21_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_22_nl = MUX_v_32_2_2(out_tmp_value_13_31_0_lpi_1_dfm_10,
      out_tmp_value_4_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_4_31_0_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_22_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_23_nl = MUX_v_32_2_2(out_tmp_value_13_31_0_lpi_1_dfm_11,
      out_tmp_value_4_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_4_63_32_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_23_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_24_nl = MUX_v_32_2_2(out_tmp_value_12_63_32_lpi_1_dfm_10,
      out_tmp_value_3_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_3_31_0_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_24_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_25_nl = MUX_v_32_2_2(out_tmp_value_12_63_32_lpi_1_dfm_11,
      out_tmp_value_3_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_3_63_32_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_25_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_26_nl = MUX_v_32_2_2(out_tmp_value_12_31_0_lpi_1_dfm_10,
      out_tmp_value_2_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_2_31_0_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_26_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_27_nl = MUX_v_32_2_2(out_tmp_value_12_31_0_lpi_1_dfm_11,
      out_tmp_value_2_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_2_63_32_lpi_1_dfm = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_27_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_28_nl = MUX_v_32_2_2(out_tmp_value_0_63_32_lpi_1_dfm_10,
      out_tmp_value_1_31_0_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_1_31_0_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_28_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_29_nl = MUX_v_32_2_2(out_tmp_value_0_63_32_lpi_1_dfm_11,
      out_tmp_value_1_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_1_63_32_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_29_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_30_nl = MUX_v_32_2_2(out_tmp_value_0_31_0_lpi_2, out_tmp_value_0_31_0_lpi_1_mx0w0,
      main_stage_0_4);
  assign out_tmp_value_0_31_0_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_30_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign out_tmp_value_mux_31_nl = MUX_v_32_2_2(out_tmp_value_0_31_0_lpi_1_dfm_10,
      out_tmp_value_0_63_32_lpi_1_mx0w0, main_stage_0_4);
  assign out_tmp_value_0_63_32_lpi_1_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      (out_tmp_value_mux_31_nl), lfst_exit_for_for_1_lpi_1_dfm_4);
  assign for_for_for_1_and_10_m1c = unequal_tmp_7 & for_for_for_1_nor_dfs_7;
  assign pe_y_reg_value_15_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_15_63_32_lpi_1_dfm_mx0,
      ({{16{COL_16_COMP_tmp_acc_psp_sva[15]}}, COL_16_COMP_tmp_acc_psp_sva}), COMP_i_0_lpi_1_dfm_6);
  assign pe_y_reg_value_15_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_16_COMP_tmp_acc_psp_sva[15]}},
      COL_16_COMP_tmp_acc_psp_sva}), pe_y_reg_value_15_31_0_lpi_1_dfm_mx0, COMP_i_0_lpi_1_dfm_6);
  assign pe_y_reg_value_14_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_14_63_32_lpi_1_dfm_mx0,
      ({{16{COL_15_COMP_tmp_acc_psp_sva[15]}}, COL_15_COMP_tmp_acc_psp_sva}), COMP_i_0_15_lpi_1_dfm_6);
  assign pe_y_reg_value_14_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_15_COMP_tmp_acc_psp_sva[15]}},
      COL_15_COMP_tmp_acc_psp_sva}), pe_y_reg_value_14_31_0_lpi_1_dfm_mx0, COMP_i_0_15_lpi_1_dfm_6);
  assign pe_y_reg_value_13_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_13_63_32_lpi_1_dfm_mx0,
      ({{16{COL_14_COMP_tmp_acc_psp_sva[15]}}, COL_14_COMP_tmp_acc_psp_sva}), COMP_i_0_14_lpi_1_dfm_6);
  assign pe_y_reg_value_13_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_14_COMP_tmp_acc_psp_sva[15]}},
      COL_14_COMP_tmp_acc_psp_sva}), pe_y_reg_value_13_31_0_lpi_1_dfm_mx0, COMP_i_0_14_lpi_1_dfm_6);
  assign pe_y_reg_value_12_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_12_63_32_lpi_1_dfm_mx0,
      ({{16{COL_13_COMP_tmp_acc_psp_sva[15]}}, COL_13_COMP_tmp_acc_psp_sva}), COMP_i_0_13_lpi_1_dfm_6);
  assign pe_y_reg_value_12_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_13_COMP_tmp_acc_psp_sva[15]}},
      COL_13_COMP_tmp_acc_psp_sva}), pe_y_reg_value_12_31_0_lpi_1_dfm_mx0, COMP_i_0_13_lpi_1_dfm_6);
  assign pe_y_reg_value_11_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_11_63_32_lpi_1_dfm_mx0,
      ({{16{COL_12_COMP_tmp_acc_psp_sva[15]}}, COL_12_COMP_tmp_acc_psp_sva}), COMP_i_0_12_lpi_1_dfm_6);
  assign pe_y_reg_value_11_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_12_COMP_tmp_acc_psp_sva[15]}},
      COL_12_COMP_tmp_acc_psp_sva}), pe_y_reg_value_11_31_0_lpi_1_dfm_mx0, COMP_i_0_12_lpi_1_dfm_6);
  assign pe_y_reg_value_10_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_10_63_32_lpi_1_dfm_mx0,
      ({{16{COL_11_COMP_tmp_acc_psp_sva[15]}}, COL_11_COMP_tmp_acc_psp_sva}), COMP_i_0_11_lpi_1_dfm_6);
  assign pe_y_reg_value_10_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_11_COMP_tmp_acc_psp_sva[15]}},
      COL_11_COMP_tmp_acc_psp_sva}), pe_y_reg_value_10_31_0_lpi_1_dfm_mx0, COMP_i_0_11_lpi_1_dfm_6);
  assign pe_y_reg_value_9_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_9_63_32_lpi_1_dfm_mx0,
      ({{16{COL_10_COMP_tmp_acc_psp_sva[15]}}, COL_10_COMP_tmp_acc_psp_sva}), COMP_i_0_10_lpi_1_dfm_6);
  assign pe_y_reg_value_9_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_10_COMP_tmp_acc_psp_sva[15]}},
      COL_10_COMP_tmp_acc_psp_sva}), pe_y_reg_value_9_31_0_lpi_1_dfm_mx0, COMP_i_0_10_lpi_1_dfm_6);
  assign pe_y_reg_value_8_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_8_63_32_lpi_1_dfm_mx0,
      ({{16{COL_9_COMP_tmp_acc_psp_sva[15]}}, COL_9_COMP_tmp_acc_psp_sva}), COMP_i_0_9_lpi_1_dfm_6);
  assign pe_y_reg_value_8_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_9_COMP_tmp_acc_psp_sva[15]}},
      COL_9_COMP_tmp_acc_psp_sva}), pe_y_reg_value_8_31_0_lpi_1_dfm_mx0, COMP_i_0_9_lpi_1_dfm_6);
  assign pe_y_reg_value_7_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_7_63_32_lpi_1_dfm_mx0,
      ({{16{COL_8_COMP_tmp_acc_psp_sva[15]}}, COL_8_COMP_tmp_acc_psp_sva}), COMP_i_0_8_lpi_1_dfm_6);
  assign pe_y_reg_value_7_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_8_COMP_tmp_acc_psp_sva[15]}},
      COL_8_COMP_tmp_acc_psp_sva}), pe_y_reg_value_7_31_0_lpi_1_dfm_mx0, COMP_i_0_8_lpi_1_dfm_6);
  assign pe_y_reg_value_6_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_6_63_32_lpi_1_dfm_mx0,
      ({{16{COL_7_COMP_tmp_acc_psp_sva[15]}}, COL_7_COMP_tmp_acc_psp_sva}), COMP_i_0_7_lpi_1_dfm_6);
  assign pe_y_reg_value_6_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_7_COMP_tmp_acc_psp_sva[15]}},
      COL_7_COMP_tmp_acc_psp_sva}), pe_y_reg_value_6_31_0_lpi_1_dfm_mx0, COMP_i_0_7_lpi_1_dfm_6);
  assign pe_y_reg_value_5_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_5_63_32_lpi_1_dfm_mx0,
      ({{16{COL_6_COMP_tmp_acc_psp_sva[15]}}, COL_6_COMP_tmp_acc_psp_sva}), COMP_i_0_6_lpi_1_dfm_6);
  assign pe_y_reg_value_5_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_6_COMP_tmp_acc_psp_sva[15]}},
      COL_6_COMP_tmp_acc_psp_sva}), pe_y_reg_value_5_31_0_lpi_1_dfm_mx0, COMP_i_0_6_lpi_1_dfm_6);
  assign pe_y_reg_value_4_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_4_63_32_lpi_1_dfm_mx0,
      ({{16{COL_5_COMP_tmp_acc_psp_sva[15]}}, COL_5_COMP_tmp_acc_psp_sva}), COMP_i_0_5_lpi_1_dfm_6);
  assign pe_y_reg_value_4_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_5_COMP_tmp_acc_psp_sva[15]}},
      COL_5_COMP_tmp_acc_psp_sva}), pe_y_reg_value_4_31_0_lpi_1_dfm_mx0, COMP_i_0_5_lpi_1_dfm_6);
  assign pe_y_reg_value_3_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_3_63_32_lpi_1_dfm_mx0,
      ({{16{COL_4_COMP_tmp_acc_psp_sva[15]}}, COL_4_COMP_tmp_acc_psp_sva}), COMP_i_0_4_lpi_1_dfm_6);
  assign pe_y_reg_value_3_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_4_COMP_tmp_acc_psp_sva[15]}},
      COL_4_COMP_tmp_acc_psp_sva}), pe_y_reg_value_3_31_0_lpi_1_dfm_mx0, COMP_i_0_4_lpi_1_dfm_6);
  assign pe_y_reg_value_2_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_2_63_32_lpi_1_dfm_mx0,
      ({{16{COL_3_COMP_tmp_acc_psp_sva[15]}}, COL_3_COMP_tmp_acc_psp_sva}), COMP_i_0_3_lpi_1_dfm_6);
  assign pe_y_reg_value_2_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_3_COMP_tmp_acc_psp_sva[15]}},
      COL_3_COMP_tmp_acc_psp_sva}), pe_y_reg_value_2_31_0_lpi_1_dfm_mx0, COMP_i_0_3_lpi_1_dfm_6);
  assign pe_y_reg_value_1_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_1_63_32_lpi_1_dfm_mx0,
      ({{16{COL_2_COMP_tmp_acc_psp_sva[15]}}, COL_2_COMP_tmp_acc_psp_sva}), COMP_i_0_2_lpi_1_dfm_6);
  assign pe_y_reg_value_1_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_2_COMP_tmp_acc_psp_sva[15]}},
      COL_2_COMP_tmp_acc_psp_sva}), pe_y_reg_value_1_31_0_lpi_1_dfm_mx0, COMP_i_0_2_lpi_1_dfm_6);
  assign pe_y_reg_value_0_63_32_sva_1_mx0 = MUX_v_32_2_2(pe_y_reg_value_0_63_32_lpi_1_dfm_mx0,
      ({{16{COL_1_COMP_tmp_acc_psp_sva[15]}}, COL_1_COMP_tmp_acc_psp_sva}), COMP_i_0_1_lpi_1_dfm_6);
  assign pe_y_reg_value_0_31_0_sva_1_mx0 = MUX_v_32_2_2(({{16{COL_1_COMP_tmp_acc_psp_sva[15]}},
      COL_1_COMP_tmp_acc_psp_sva}), pe_y_reg_value_0_31_0_lpi_1_dfm_mx0, COMP_i_0_1_lpi_1_dfm_6);
  assign pe_y_reg_value_15_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_15_63_32_lpi_2,
      out_tmp_value_15_63_32_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_16_COMP_tmp_mul_nl = $signed(in_tmp_16_lpi_1_dfm_5) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_16_COMP_tmp_mul_nl = nl_COL_16_COMP_tmp_mul_nl[15:0];
  assign nl_COL_16_COMP_tmp_acc_psp_sva = (COL_16_COMP_tmp_mul_nl) + COL_16_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_16_COMP_tmp_acc_psp_sva = nl_COL_16_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_15_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_15_31_0_lpi_2,
      out_tmp_value_15_31_0_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign in_tmp_16_lpi_1_dfm_1 = MUX1HOT_v_16_3_2(in_tmp_16_lpi_2, (input_rsci_d_mxwt[255:240]),
      (input_rsci_d_mxwt[15:0]), {(~ exitL_exit_COL_1_COMP_lpi_1_dfm_4) , asn_259
      , asn_261});
  assign pe_y_reg_value_14_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_14_63_32_lpi_2,
      out_tmp_value_14_63_32_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_15_COMP_tmp_mul_nl = $signed(mux_63_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_15_COMP_tmp_mul_nl = nl_COL_15_COMP_tmp_mul_nl[15:0];
  assign nl_COL_15_COMP_tmp_acc_psp_sva = (COL_15_COMP_tmp_mul_nl) + COL_15_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_15_COMP_tmp_acc_psp_sva = nl_COL_15_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_14_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_14_31_0_lpi_2,
      out_tmp_value_14_31_0_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_13_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_13_63_32_lpi_2,
      out_tmp_value_13_63_32_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_14_COMP_tmp_mul_nl = $signed(mux_48_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_14_COMP_tmp_mul_nl = nl_COL_14_COMP_tmp_mul_nl[15:0];
  assign nl_COL_14_COMP_tmp_acc_psp_sva = (COL_14_COMP_tmp_mul_nl) + COL_14_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_14_COMP_tmp_acc_psp_sva = nl_COL_14_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_13_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_13_31_0_lpi_2,
      out_tmp_value_13_31_0_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_12_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_12_63_32_lpi_2,
      out_tmp_value_12_63_32_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_13_COMP_tmp_mul_nl = $signed(mux_47_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_13_COMP_tmp_mul_nl = nl_COL_13_COMP_tmp_mul_nl[15:0];
  assign nl_COL_13_COMP_tmp_acc_psp_sva = (COL_13_COMP_tmp_mul_nl) + COL_13_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_13_COMP_tmp_acc_psp_sva = nl_COL_13_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_12_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_12_31_0_lpi_2,
      out_tmp_value_12_31_0_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_11_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_11_63_32_lpi_2,
      out_tmp_value_11_63_32_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_12_COMP_tmp_mul_nl = $signed(mux_46_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_12_COMP_tmp_mul_nl = nl_COL_12_COMP_tmp_mul_nl[15:0];
  assign nl_COL_12_COMP_tmp_acc_psp_sva = (COL_12_COMP_tmp_mul_nl) + COL_12_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_12_COMP_tmp_acc_psp_sva = nl_COL_12_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_11_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_11_31_0_lpi_2,
      out_tmp_value_11_31_0_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_10_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_10_63_32_lpi_2,
      out_tmp_value_10_63_32_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_11_COMP_tmp_mul_nl = $signed(mux_45_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_11_COMP_tmp_mul_nl = nl_COL_11_COMP_tmp_mul_nl[15:0];
  assign nl_COL_11_COMP_tmp_acc_psp_sva = (COL_11_COMP_tmp_mul_nl) + COL_11_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_11_COMP_tmp_acc_psp_sva = nl_COL_11_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_10_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_10_31_0_lpi_2,
      out_tmp_value_10_31_0_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_9_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_9_63_32_lpi_2,
      out_tmp_value_9_63_32_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_10_COMP_tmp_mul_nl = $signed(mux_44_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_10_COMP_tmp_mul_nl = nl_COL_10_COMP_tmp_mul_nl[15:0];
  assign nl_COL_10_COMP_tmp_acc_psp_sva = (COL_10_COMP_tmp_mul_nl) + COL_10_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_10_COMP_tmp_acc_psp_sva = nl_COL_10_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_9_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_9_31_0_lpi_2,
      out_tmp_value_9_31_0_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_8_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_8_63_32_lpi_2,
      out_tmp_value_8_63_32_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_9_COMP_tmp_mul_nl = $signed(mux_43_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_9_COMP_tmp_mul_nl = nl_COL_9_COMP_tmp_mul_nl[15:0];
  assign nl_COL_9_COMP_tmp_acc_psp_sva = (COL_9_COMP_tmp_mul_nl) + COL_9_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_9_COMP_tmp_acc_psp_sva = nl_COL_9_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_8_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_8_31_0_lpi_2,
      out_tmp_value_8_31_0_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_7_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_7_63_32_lpi_2,
      out_tmp_value_7_63_32_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_8_COMP_tmp_mul_nl = $signed(mux_42_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_8_COMP_tmp_mul_nl = nl_COL_8_COMP_tmp_mul_nl[15:0];
  assign nl_COL_8_COMP_tmp_acc_psp_sva = (COL_8_COMP_tmp_mul_nl) + COL_8_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_8_COMP_tmp_acc_psp_sva = nl_COL_8_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_7_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_7_31_0_lpi_2,
      out_tmp_value_7_31_0_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_6_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_6_63_32_lpi_2,
      out_tmp_value_6_63_32_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_7_COMP_tmp_mul_nl = $signed(mux_41_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_7_COMP_tmp_mul_nl = nl_COL_7_COMP_tmp_mul_nl[15:0];
  assign nl_COL_7_COMP_tmp_acc_psp_sva = (COL_7_COMP_tmp_mul_nl) + COL_7_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_7_COMP_tmp_acc_psp_sva = nl_COL_7_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_6_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_6_31_0_lpi_2,
      out_tmp_value_6_31_0_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_5_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_5_63_32_lpi_2,
      out_tmp_value_5_63_32_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_6_COMP_tmp_mul_nl = $signed(mux_40_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_6_COMP_tmp_mul_nl = nl_COL_6_COMP_tmp_mul_nl[15:0];
  assign nl_COL_6_COMP_tmp_acc_psp_sva = (COL_6_COMP_tmp_mul_nl) + COL_6_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_6_COMP_tmp_acc_psp_sva = nl_COL_6_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_5_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_5_31_0_lpi_2,
      out_tmp_value_5_31_0_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_4_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_4_63_32_lpi_2,
      out_tmp_value_4_63_32_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_5_COMP_tmp_mul_nl = $signed(mux_39_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_5_COMP_tmp_mul_nl = nl_COL_5_COMP_tmp_mul_nl[15:0];
  assign nl_COL_5_COMP_tmp_acc_psp_sva = (COL_5_COMP_tmp_mul_nl) + COL_5_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_5_COMP_tmp_acc_psp_sva = nl_COL_5_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_4_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_4_31_0_lpi_2,
      out_tmp_value_4_31_0_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_3_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_3_63_32_lpi_2,
      out_tmp_value_3_63_32_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_4_COMP_tmp_mul_nl = $signed(mux_38_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_4_COMP_tmp_mul_nl = nl_COL_4_COMP_tmp_mul_nl[15:0];
  assign nl_COL_4_COMP_tmp_acc_psp_sva = (COL_4_COMP_tmp_mul_nl) + COL_4_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_4_COMP_tmp_acc_psp_sva = nl_COL_4_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_3_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_3_31_0_lpi_2,
      out_tmp_value_3_31_0_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_2_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_2_63_32_lpi_2,
      out_tmp_value_2_63_32_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_3_COMP_tmp_mul_nl = $signed(mux_37_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_3_COMP_tmp_mul_nl = nl_COL_3_COMP_tmp_mul_nl[15:0];
  assign nl_COL_3_COMP_tmp_acc_psp_sva = (COL_3_COMP_tmp_mul_nl) + COL_3_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_3_COMP_tmp_acc_psp_sva = nl_COL_3_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_2_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_2_31_0_lpi_2,
      out_tmp_value_2_31_0_lpi_1_dfm, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_1_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_1_63_32_lpi_2,
      out_tmp_value_1_63_32_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_2_COMP_tmp_mul_nl = $signed(mux_36_itm_2) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_2_COMP_tmp_mul_nl = nl_COL_2_COMP_tmp_mul_nl[15:0];
  assign nl_COL_2_COMP_tmp_acc_psp_sva = (COL_2_COMP_tmp_mul_nl) + COL_2_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_2_COMP_tmp_acc_psp_sva = nl_COL_2_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_1_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_1_31_0_lpi_2,
      out_tmp_value_1_31_0_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_y_reg_value_0_63_32_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_0_63_32_lpi_2,
      out_tmp_value_0_63_32_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign nl_COL_1_COMP_tmp_mul_nl = $signed(pe_x_reg_0_lpi_1_dfm_4) * $signed(conv_u2s_16_17(COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000));
  assign COL_1_COMP_tmp_mul_nl = nl_COL_1_COMP_tmp_mul_nl[15:0];
  assign nl_COL_1_COMP_tmp_acc_psp_sva = (COL_1_COMP_tmp_mul_nl) + COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_2_rshift_itm;
  assign COL_1_COMP_tmp_acc_psp_sva = nl_COL_1_COMP_tmp_acc_psp_sva[15:0];
  assign pe_y_reg_value_0_31_0_lpi_1_dfm_mx0 = MUX_v_32_2_2(pe_y_reg_value_0_31_0_lpi_2,
      out_tmp_value_0_31_0_lpi_1_dfm_mx0w0, exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign pe_x_reg_0_lpi_1_dfm = MUX1HOT_v_16_3_2(pe_x_reg_0_lpi_2, (input_rsci_d_mxwt[15:0]),
      in_tmp_1_lpi_2, {(~ exitL_exit_COL_1_COMP_lpi_1_dfm_4) , asn_259 , asn_261});
  assign unequal_tmp = (WY_mux_3_cse!=2'b00);
  assign nl_for_acc_2_tmp = conv_u2u_2_3(for_ko_2_0_lpi_1_dfm_1_0) + 3'b1;
  assign for_acc_2_tmp = nl_for_acc_2_tmp[2:0];
  assign for_for_for_1_equal_tmp = lfst_exit_for_for_for_1_lpi_1_dfm_1 & (~ lfst_exit_for_for_for_1_lpi_1_dfm_0);
  assign for_for_for_1_and_4_m1c = unequal_tmp & for_for_for_1_nor_dfs;
  assign for_for_for_1_equal_tmp_1 = lfst_exit_for_for_for_1_lpi_1_dfm_1 & lfst_exit_for_for_for_1_lpi_1_dfm_0;
  assign for_for_for_1_and_3_cse = (~ unequal_tmp) & for_for_for_1_nor_dfs;
  assign for_for_for_1_and_96_cse = (~ exit_for_for_for_1_lpi_1_dfm_1) & for_for_for_1_equal_tmp;
  assign for_for_for_1_and_95_cse = exit_for_for_for_1_lpi_1_dfm_1 & for_for_for_1_equal_tmp;
  assign for_for_for_1_and_2_m1c = (~ exit_for_for_lpi_1_dfm_5) & for_for_for_1_equal_tmp;
  assign for_for_for_1_nor_dfs = ~(for_for_for_1_equal_tmp | for_for_for_1_equal_tmp_1);
  assign for_for_for_1_and_97_cse = for_for_for_1_for_q_0_lpi_2 & for_for_for_1_equal_tmp;
  assign for_not_39_nl = ~ exitL_exit_for_sva;
  assign for_ko_2_0_lpi_1_dfm_1_0 = MUX_v_2_2_2(2'b00, for_ko_2_0_lpi_1_1_0_1, (for_not_39_nl));
  assign WX_and_16_psp_mx0w0 = WX_if_1_and_stg_2_0_sva_mx0 & (WX_if_1_acc_decb_sva_1_3_1_1[2])
      & (~ WX_unequal_tmp_1);
  assign WX_and_14_psp_mx0w0 = WX_if_1_and_stg_1_3_sva_mx0 & (WX_if_1_acc_decb_sva_1_3_1_1[2:1]==2'b01)
      & (~ WX_unequal_tmp_1);
  assign WX_and_12_psp_mx0w0 = WX_if_1_and_stg_1_2_sva_mx0 & (WX_if_1_acc_decb_sva_1_3_1_1[2:1]==2'b01)
      & (~ WX_unequal_tmp_1);
  assign WX_and_10_psp_mx0w0 = WX_if_1_and_stg_1_1_sva_mx0 & (WX_if_1_acc_decb_sva_1_3_1_1[2:1]==2'b01)
      & (~ WX_unequal_tmp_1);
  assign WX_if_1_mux_26_nl = MUX_s_1_2_2(WX_if_1_and_stg_1_0_sva_mx0w0, WX_if_1_and_stg_1_0_sva,
      or_dcpl_76);
  assign WX_and_8_psp_mx0w0 = (WX_if_1_mux_26_nl) & (WX_if_1_acc_decb_sva_1_3_1_1[2:1]==2'b01)
      & (~ WX_unequal_tmp_1);
  assign WX_and_6_psp_mx0w0 = ~((~ WX_if_1_and_stg_1_3_sva_mx0) | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b00)
      | WX_unequal_tmp_1);
  assign WX_and_4_psp_mx0w0 = ~((~ WX_if_1_and_stg_1_2_sva_mx0) | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b00)
      | WX_unequal_tmp_1);
  assign WX_and_2_psp_mx0w0 = ~((~ WX_if_1_and_stg_1_1_sva_mx0) | (WX_if_1_acc_decb_sva_1_3_1_1[2:1]!=2'b00)
      | WX_unequal_tmp_1);
  assign WX_and_psp_mx0w0 = WX_if_1_and_stg_2_0_sva_mx0 & (~ (WX_if_1_acc_decb_sva_1_3_1_1[2]))
      & (~ WX_unequal_tmp_1);
  assign in_tmp_14_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[223:208]), in_tmp_14_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_13_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[207:192]), in_tmp_13_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_12_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[191:176]), in_tmp_12_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_11_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[175:160]), in_tmp_11_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_10_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[159:144]), in_tmp_10_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_9_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[143:128]), in_tmp_9_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_8_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[127:112]), in_tmp_8_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_7_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[111:96]), in_tmp_7_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_6_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[95:80]), in_tmp_6_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_5_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[79:64]), in_tmp_5_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_4_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[63:48]), in_tmp_4_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_3_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[47:32]), in_tmp_3_lpi_2,
      WX_unequal_tmp_5);
  assign in_tmp_2_lpi_1_dfm_1_mx0 = MUX_v_16_2_2((input_rsci_d_mxwt[31:16]), in_tmp_2_lpi_2,
      WX_unequal_tmp_5);
  assign WX_if_1_and_stg_1_1_sva_mx0w0 = out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1
      & (~ (WX_if_1_acc_decb_sva_1_3_1_1[0]));
  assign WX_if_1_and_stg_1_1_sva_mx0 = MUX_s_1_2_2(WX_if_1_and_stg_1_1_sva_mx0w0,
      WX_if_1_and_stg_1_1_sva, or_dcpl_76);
  assign WX_if_1_and_stg_1_2_sva_mx0w0 = (~ out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1)
      & (WX_if_1_acc_decb_sva_1_3_1_1[0]);
  assign WX_if_1_and_stg_1_2_sva_mx0 = MUX_s_1_2_2(WX_if_1_and_stg_1_2_sva_mx0w0,
      WX_if_1_and_stg_1_2_sva, or_dcpl_76);
  assign WX_if_1_and_stg_1_3_sva_mx0w0 = out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1
      & (WX_if_1_acc_decb_sva_1_3_1_1[0]);
  assign WX_if_1_and_stg_1_3_sva_mx0 = MUX_s_1_2_2(WX_if_1_and_stg_1_3_sva_mx0w0,
      WX_if_1_and_stg_1_3_sva, or_dcpl_76);
  assign WX_if_1_and_stg_2_0_sva_mx0w0 = WX_if_1_and_stg_1_0_sva_mx0w0 & (~ (WX_if_1_acc_decb_sva_1_3_1_1[1]));
  assign WX_if_1_and_stg_2_0_sva_mx0 = MUX_s_1_2_2(WX_if_1_and_stg_2_0_sva_mx0w0,
      WX_if_1_and_stg_2_0_sva, or_dcpl_76);
  assign WX_if_1_and_stg_1_0_sva_mx0w0 = ~(out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1
      | (WX_if_1_acc_decb_sva_1_3_1_1[0]));
  assign nl_WX_if_1_acc_decb_sva_3_1_mx0w0 = conv_u2u_2_3(WX_if_1_acc_1_ncse[2:1])
      + conv_u2u_2_3(WY_wy_1_0_lpi_1_dfm);
  assign WX_if_1_acc_decb_sva_3_1_mx0w0 = nl_WX_if_1_acc_decb_sva_3_1_mx0w0[2:0];
  assign WX_unequal_tmp_1 = (for_for_row_6_0_lpi_1_dfm_9[5:0]!=6'b000000);
  assign asn_259 = (~ WX_unequal_tmp_5) & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign for_for_for_1_or_cse = for_for_for_1_equal_tmp_2 | for_for_for_1_equal_tmp_5;
  assign nl_WX_if_1_acc_1_ncse = conv_u2u_2_3(WY_wy_1_0_lpi_1_dfm) + conv_u2u_2_3(WX_wx_1_0_lpi_1_dfm);
  assign WX_if_1_acc_1_ncse = nl_WX_if_1_acc_1_ncse[2:0];
  assign for_for_for_1_asn_426 = (~ unequal_tmp_7) & for_for_for_1_nor_dfs_7;
  assign for_for_for_1_asn_428 = ((~ COMP_and_13_mdf_sva_7) & for_for_for_1_and_10_m1c)
      | (lfst_exit_for_for_for_1_lpi_1_dfm_10_1_1 & for_for_for_1_equal_tmp_11) |
      for_for_for_1_equal_tmp_13;
  assign for_for_for_1_asn_430 = COMP_and_13_mdf_sva_7 & for_for_for_1_and_10_m1c;
  assign for_for_for_1_asn_432 = (~ lfst_exit_for_for_for_1_lpi_1_dfm_10_1_1) & for_for_for_1_equal_tmp_11;
  assign asn_261 = WX_unequal_tmp_5 & exitL_exit_COL_1_COMP_lpi_1_dfm_4;
  assign WY_mux_6_tmp = MUX_v_2_2_2(2'b1, 2'b10, exit_WY_lpi_1_dfm_2);
  assign and_dcpl_1 = (~ lfst_exit_for_for_for_1_lpi_1_dfm_st_1_0) & lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1;
  assign or_dcpl = ~(main_stage_0_2 & for_for_for_1_equal_tmp_2);
  assign or_tmp_4 = nor_41_cse | (~ lfst_exit_for_for_1_lpi_2) | exitL_exit_for_sva
      | exit_for_lpi_1_dfm_4;
  assign or_tmp_5 = main_stage_0_2 | (~ or_tmp_4);
  assign mux_tmp = MUX_s_1_2_2((~ or_tmp_4), for_for_for_1_equal_tmp_5, main_stage_0_2);
  assign or_dcpl_7 = exit_for_lpi_1_dfm_4 | exitL_exit_for_sva;
  assign or_dcpl_9 = ~((for_for_acc_1_tmp[6]) & (for_acc_2_tmp[2]));
  assign or_dcpl_13 = or_dcpl_7 | (~ lfst_exit_for_for_1_lpi_2);
  assign or_dcpl_14 = or_dcpl_13 | (~ lfst_exit_for_for_for_1_lpi_1_1_1) | lfst_exit_for_for_for_1_lpi_1_0_1;
  assign or_dcpl_15 = or_dcpl_14 | (~((for_for_for_1_acc_1_tmp[4]) & for_for_for_1_for_q_0_lpi_2))
      | or_dcpl_9;
  assign nor_53_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1);
  assign mux_153_nl = MUX_s_1_2_2((nor_53_nl), COMP_and_13_mdf_sva_6, unequal_tmp_6);
  assign and_dcpl_15 = (mux_153_nl) & or_395_cse & for_for_for_1_nor_dfs_6 & main_stage_0_3;
  assign and_dcpl_27 = (~ or_dcpl_13) & lfst_exit_for_for_for_1_lpi_1_1_1 & (~ lfst_exit_for_for_for_1_lpi_1_0_1);
  assign or_dcpl_18 = or_dcpl_13 | (~ lfst_exit_for_for_for_1_lpi_1_1_1) | (~ lfst_exit_for_for_for_1_lpi_1_0_1);
  assign and_dcpl_36 = (~ lfst_exit_for_for_for_1_lpi_1_1_1) & lfst_exit_for_for_for_1_lpi_1_0_1;
  assign or_tmp_16 = (~ lfst_exit_WX_1_lpi_1) | exitL_exit_COL_1_COMP_lpi_1;
  assign and_tmp_2 = ((WX_wx_1_0_lpi_3!=2'b00)) & or_tmp_16;
  assign or_tmp_19 = (WX_wx_1_0_lpi_3!=2'b00) | (~ or_tmp_16);
  assign or_41_nl = (~ COMP_and_13_tmp) | (for_for_for_1_for_for_for_1_for_for_for_1_mux1h_1_tmp!=2'b00);
  assign mux_157_nl = MUX_s_1_2_2(and_tmp_2, or_tmp_19, or_41_nl);
  assign or_38_nl = (~ for_for_for_1_nand_2_tmp) | (WY_mux_6_tmp!=2'b01);
  assign mux_158_nl = MUX_s_1_2_2((mux_157_nl), and_tmp_2, or_38_nl);
  assign and_dcpl_38 = (mux_158_nl) & (~ or_dcpl_13) & and_dcpl_36;
  assign and_dcpl_48 = lfst_exit_for_lpi_1_dfm & lfst_exit_for_for_1_lpi_2 & (~ lfst_exit_for_for_for_1_lpi_1_1_1)
      & lfst_exit_for_for_for_1_lpi_1_0_1 & (~ exitL_exit_COL_1_COMP_lpi_1) & lfst_exit_WX_1_lpi_1;
  assign or_dcpl_28 = (~(lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 & main_stage_0_3))
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_0_1 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4);
  assign and_dcpl_59 = lfst_exit_for_for_for_1_lpi_1_0_1 & (~ exitL_exit_COL_1_COMP_lpi_1)
      & lfst_exit_WX_1_lpi_1;
  assign or_dcpl_35 = and_dcpl_59 | lfst_exit_for_for_for_1_lpi_1_1_1;
  assign and_dcpl_61 = ((or_dcpl_35 & lfst_exit_for_for_1_lpi_2) | (for_for_row_6_0_lpi_3[5:0]!=6'b000000))
      & lfst_exit_for_lpi_1_dfm;
  assign and_dcpl_63 = or_dcpl_35 & lfst_exit_for_for_1_lpi_1_dfm;
  assign or_dcpl_38 = (~ COMP_and_13_tmp) | WX_acc_tmp_1;
  assign and_dcpl_65 = lfst_exit_for_lpi_1_dfm & lfst_exit_for_for_1_lpi_2 & lfst_exit_for_for_for_1_lpi_1_1_1;
  assign and_dcpl_66 = (~ main_stage_0_3) & main_stage_0_4;
  assign and_dcpl_68 = COMP_and_13_mdf_sva_6 & (~ unequal_tmp_6);
  assign and_dcpl_69 = COMP_and_13_mdf_sva_6 & unequal_tmp_6;
  assign and_dcpl_70 = and_dcpl_69 & COMP_i_0_7_lpi_1_dfm_6;
  assign and_dcpl_71 = and_dcpl_69 & (~ COMP_i_0_7_lpi_1_dfm_6);
  assign and_dcpl_72 = and_dcpl_69 & COMP_i_0_6_lpi_1_dfm_6;
  assign and_dcpl_73 = and_dcpl_69 & (~ COMP_i_0_6_lpi_1_dfm_6);
  assign and_dcpl_74 = and_dcpl_69 & COMP_i_0_5_lpi_1_dfm_6;
  assign and_dcpl_75 = and_dcpl_69 & (~ COMP_i_0_5_lpi_1_dfm_6);
  assign and_dcpl_76 = and_dcpl_69 & COMP_i_0_4_lpi_1_dfm_6;
  assign and_dcpl_77 = and_dcpl_69 & (~ COMP_i_0_4_lpi_1_dfm_6);
  assign and_dcpl_78 = and_dcpl_69 & COMP_i_0_3_lpi_1_dfm_6;
  assign and_dcpl_79 = and_dcpl_69 & (~ COMP_i_0_3_lpi_1_dfm_6);
  assign and_dcpl_80 = and_dcpl_69 & COMP_i_0_lpi_1_dfm_6;
  assign and_dcpl_81 = and_dcpl_69 & (~ COMP_i_0_lpi_1_dfm_6);
  assign and_dcpl_82 = and_dcpl_69 & COMP_i_0_15_lpi_1_dfm_6;
  assign and_dcpl_83 = and_dcpl_69 & (~ COMP_i_0_15_lpi_1_dfm_6);
  assign and_dcpl_84 = and_dcpl_69 & COMP_i_0_14_lpi_1_dfm_6;
  assign and_dcpl_85 = and_dcpl_69 & (~ COMP_i_0_14_lpi_1_dfm_6);
  assign and_dcpl_86 = and_dcpl_69 & COMP_i_0_13_lpi_1_dfm_6;
  assign and_dcpl_87 = and_dcpl_69 & (~ COMP_i_0_13_lpi_1_dfm_6);
  assign and_dcpl_88 = and_dcpl_69 & COMP_i_0_12_lpi_1_dfm_6;
  assign and_dcpl_89 = and_dcpl_69 & (~ COMP_i_0_12_lpi_1_dfm_6);
  assign and_dcpl_90 = and_dcpl_69 & COMP_i_0_11_lpi_1_dfm_6;
  assign and_dcpl_91 = and_dcpl_69 & (~ COMP_i_0_11_lpi_1_dfm_6);
  assign and_dcpl_92 = and_dcpl_69 & COMP_i_0_2_lpi_1_dfm_6;
  assign and_dcpl_93 = and_dcpl_69 & (~ COMP_i_0_2_lpi_1_dfm_6);
  assign and_dcpl_94 = and_dcpl_69 & COMP_i_0_1_lpi_1_dfm_6;
  assign and_dcpl_95 = and_dcpl_69 & (~ COMP_i_0_1_lpi_1_dfm_6);
  assign and_dcpl_96 = and_dcpl_69 & COMP_i_0_10_lpi_1_dfm_6;
  assign and_dcpl_97 = and_dcpl_69 & (~ COMP_i_0_10_lpi_1_dfm_6);
  assign and_dcpl_98 = and_dcpl_69 & COMP_i_0_9_lpi_1_dfm_6;
  assign and_dcpl_99 = and_dcpl_69 & (~ COMP_i_0_9_lpi_1_dfm_6);
  assign and_dcpl_100 = and_dcpl_69 & COMP_i_0_8_lpi_1_dfm_6;
  assign and_dcpl_101 = and_dcpl_69 & (~ COMP_i_0_8_lpi_1_dfm_6);
  assign or_dcpl_50 = (~ main_stage_0_2) | for_for_for_1_equal_tmp_5;
  assign or_dcpl_51 = or_dcpl_50 | for_for_for_1_equal_tmp_2 | (~ exitL_exit_COL_1_COMP_lpi_1_dfm_4);
  assign or_dcpl_70 = ~(main_stage_0_2 & exitL_exit_COL_1_COMP_lpi_1_dfm_4);
  assign or_dcpl_72 = (for_for_row_slc_for_for_row_6_0_5_0_1_itm_3[1:0]!=2'b00);
  assign or_dcpl_76 = (for_for_row_slc_for_for_row_6_0_5_0_1_itm_3[3]) | (for_for_row_slc_for_for_row_6_0_5_0_1_itm_3[5])
      | (for_for_row_slc_for_for_row_6_0_5_0_1_itm_3[2]) | or_dcpl_72 | (for_for_row_slc_for_for_row_6_0_5_0_1_itm_3[4]);
  assign or_tmp_84 = lfst_exit_for_for_for_1_lpi_1_dfm_9_1_1 | nand_75_cse;
  assign not_tmp_131 = ~((for_for_for_1_nor_dfs_7 | for_for_for_1_equal_tmp_11 |
      for_for_for_1_equal_tmp_13) & main_stage_0_4);
  assign or_tmp_250 = (~ lfst_exit_for_for_1_lpi_1_dfm_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13 | (~ main_stage_0_4);
  assign mux_414_cse = MUX_v_16_2_2((weight_rsci_d_mxwt[15:0]), (weight_rsci_d_mxwt[31:16]),
      COMP_i_0_1_lpi_1_dfm_5);
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_1_asn_itm_2 <= {512'b0 , 512'b0};
    end
    else if ( core_wen & main_stage_0_3 & for_for_for_1_equal_tmp_10 & (or_dcpl |
        and_dcpl_1) ) begin
      for_for_for_1_asn_itm_2 <= for_for_out_stencil_value_sva_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_1_equal_tmp_11 <= 1'b0;
    end
    else if ( core_wen & (or_dcpl | lfst_exit_for_for_1_lpi_1_dfm_1 | and_dcpl_1)
        & main_stage_0_3 ) begin
      for_for_for_1_equal_tmp_11 <= for_for_for_1_equal_tmp_10;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_output_rsci_oswt_cse <= 1'b0;
      lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1 <= 1'b0;
      lfst_exit_for_for_for_1_lpi_1_dfm_st_1_0 <= 1'b0;
      reg_weight_rsci_oswt_cse <= 1'b0;
      reg_input_rsci_oswt_cse <= 1'b0;
      lfst_exit_for_for_for_1_lpi_1_1_1 <= 1'b0;
      lfst_exit_for_for_for_1_lpi_1_0_1 <= 1'b0;
      lfst_exit_for_for_1_lpi_2 <= 1'b0;
      exit_for_lpi_1_dfm_4 <= 1'b0;
      exitL_exit_for_sva <= 1'b1;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      slc_lfst_exit_for_for_for_1_1_1_itm_4 <= 1'b0;
      for_for_for_1_equal_tmp_5 <= 1'b0;
      for_for_for_1_equal_tmp_2 <= 1'b0;
      lfst_exit_for_for_1_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_output_rsci_oswt_cse <= ~ or_dcpl_28;
      lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1 <= lfst_exit_for_for_for_1_lpi_1_dfm_1;
      lfst_exit_for_for_for_1_lpi_1_dfm_st_1_0 <= lfst_exit_for_for_for_1_lpi_1_dfm_0;
      reg_weight_rsci_oswt_cse <= ~ and_dcpl_61;
      reg_input_rsci_oswt_cse <= ~ and_dcpl_63;
      lfst_exit_for_for_for_1_lpi_1_1_1 <= (for_for_for_1_mux1h_196_nl) & (~ for_for_for_1_and_95_cse);
      lfst_exit_for_for_for_1_lpi_1_0_1 <= (for_for_for_1_mux1h_193_nl) & (~(for_for_for_1_and_95_cse
          | for_for_for_1_and_96_cse));
      lfst_exit_for_for_1_lpi_2 <= for_for_for_1_nand_2_tmp;
      exit_for_lpi_1_dfm_4 <= exit_for_lpi_1_dfm_3;
      exitL_exit_for_sva <= exit_for_lpi_1_dfm_3;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      slc_lfst_exit_for_for_for_1_1_1_itm_4 <= ~ exit_for_for_for_1_lpi_1_dfm_1;
      for_for_for_1_equal_tmp_5 <= for_for_for_1_equal_tmp_1;
      for_for_for_1_equal_tmp_2 <= for_for_for_1_equal_tmp;
      lfst_exit_for_for_1_lpi_1_dfm_1 <= lfst_exit_for_for_1_lpi_1_dfm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      output_rsci_d <= {512'b0 , 512'b0};
    end
    else if ( core_wen & (~ or_dcpl_28) ) begin
      output_rsci_d <= for_for_out_stencil_value_sva_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5 <= 2'b0;
      COMP_i_0_lpi_1_dfm_6 <= 1'b0;
      in_tmp_16_lpi_1_dfm_5 <= 16'b0;
      COMP_i_0_15_lpi_1_dfm_6 <= 1'b0;
      mux_63_itm_2 <= 16'b0;
      COMP_i_0_14_lpi_1_dfm_6 <= 1'b0;
      mux_48_itm_2 <= 16'b0;
      COMP_i_0_13_lpi_1_dfm_6 <= 1'b0;
      mux_47_itm_2 <= 16'b0;
      COMP_i_0_12_lpi_1_dfm_6 <= 1'b0;
      mux_46_itm_2 <= 16'b0;
      COMP_i_0_11_lpi_1_dfm_6 <= 1'b0;
      mux_45_itm_2 <= 16'b0;
      COMP_i_0_10_lpi_1_dfm_6 <= 1'b0;
      mux_44_itm_2 <= 16'b0;
      COMP_i_0_9_lpi_1_dfm_6 <= 1'b0;
      mux_43_itm_2 <= 16'b0;
      COMP_i_0_8_lpi_1_dfm_6 <= 1'b0;
      mux_42_itm_2 <= 16'b0;
      COMP_i_0_7_lpi_1_dfm_6 <= 1'b0;
      mux_41_itm_2 <= 16'b0;
      COMP_i_0_6_lpi_1_dfm_6 <= 1'b0;
      mux_40_itm_2 <= 16'b0;
      COMP_i_0_5_lpi_1_dfm_6 <= 1'b0;
      mux_39_itm_2 <= 16'b0;
      COMP_i_0_4_lpi_1_dfm_6 <= 1'b0;
      mux_38_itm_2 <= 16'b0;
      COMP_i_0_3_lpi_1_dfm_6 <= 1'b0;
      mux_37_itm_2 <= 16'b0;
      COMP_i_0_2_lpi_1_dfm_6 <= 1'b0;
      mux_36_itm_2 <= 16'b0;
      COMP_i_0_1_lpi_1_dfm_6 <= 1'b0;
      pe_x_reg_0_lpi_1_dfm_4 <= 16'b0;
    end
    else if ( for_for_for_1_and_289_cse ) begin
      lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5 <= lfst_exit_for_for_for_1_lpi_1_dfm_1_st_4;
      COMP_i_0_lpi_1_dfm_6 <= COMP_i_0_lpi_1_dfm_5;
      in_tmp_16_lpi_1_dfm_5 <= in_tmp_16_lpi_1_dfm_1;
      COMP_i_0_15_lpi_1_dfm_6 <= COMP_i_0_15_lpi_1_dfm_5;
      mux_63_itm_2 <= MUX_v_16_2_2((input_rsci_d_mxwt[239:224]), in_tmp_15_lpi_2,
          or_68_nl);
      COMP_i_0_14_lpi_1_dfm_6 <= COMP_i_0_14_lpi_1_dfm_5;
      mux_48_itm_2 <= MUX_v_16_2_2(pe_x_reg_13_lpi_2, in_tmp_14_lpi_1_dfm_1_mx0,
          exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_13_lpi_1_dfm_6 <= COMP_i_0_13_lpi_1_dfm_5;
      mux_47_itm_2 <= MUX_v_16_2_2(pe_x_reg_12_lpi_2, in_tmp_13_lpi_1_dfm_1_mx0,
          exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_12_lpi_1_dfm_6 <= COMP_i_0_12_lpi_1_dfm_5;
      mux_46_itm_2 <= MUX_v_16_2_2(pe_x_reg_11_lpi_2, in_tmp_12_lpi_1_dfm_1_mx0,
          exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_11_lpi_1_dfm_6 <= COMP_i_0_11_lpi_1_dfm_5;
      mux_45_itm_2 <= MUX_v_16_2_2(pe_x_reg_10_lpi_2, in_tmp_11_lpi_1_dfm_1_mx0,
          exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_10_lpi_1_dfm_6 <= COMP_i_0_10_lpi_1_dfm_5;
      mux_44_itm_2 <= MUX_v_16_2_2(pe_x_reg_9_lpi_2, in_tmp_10_lpi_1_dfm_1_mx0, exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_9_lpi_1_dfm_6 <= COMP_i_0_9_lpi_1_dfm_5;
      mux_43_itm_2 <= MUX_v_16_2_2(pe_x_reg_8_lpi_2, in_tmp_9_lpi_1_dfm_1_mx0, exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_8_lpi_1_dfm_6 <= COMP_i_0_8_lpi_1_dfm_5;
      mux_42_itm_2 <= MUX_v_16_2_2(pe_x_reg_7_lpi_2, in_tmp_8_lpi_1_dfm_1_mx0, exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_7_lpi_1_dfm_6 <= COMP_i_0_7_lpi_1_dfm_5;
      mux_41_itm_2 <= MUX_v_16_2_2(pe_x_reg_6_lpi_2, in_tmp_7_lpi_1_dfm_1_mx0, exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_6_lpi_1_dfm_6 <= COMP_i_0_6_lpi_1_dfm_5;
      mux_40_itm_2 <= MUX_v_16_2_2(pe_x_reg_5_lpi_2, in_tmp_6_lpi_1_dfm_1_mx0, exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_5_lpi_1_dfm_6 <= COMP_i_0_5_lpi_1_dfm_5;
      mux_39_itm_2 <= MUX_v_16_2_2(pe_x_reg_4_lpi_2, in_tmp_5_lpi_1_dfm_1_mx0, exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_4_lpi_1_dfm_6 <= COMP_i_0_4_lpi_1_dfm_5;
      mux_38_itm_2 <= MUX_v_16_2_2(pe_x_reg_3_lpi_2, in_tmp_4_lpi_1_dfm_1_mx0, exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_3_lpi_1_dfm_6 <= COMP_i_0_3_lpi_1_dfm_5;
      mux_37_itm_2 <= MUX_v_16_2_2(pe_x_reg_2_lpi_2, in_tmp_3_lpi_1_dfm_1_mx0, exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_2_lpi_1_dfm_6 <= COMP_i_0_2_lpi_1_dfm_5;
      mux_36_itm_2 <= MUX_v_16_2_2(pe_x_reg_1_lpi_2, in_tmp_2_lpi_1_dfm_1_mx0, exitL_exit_COL_1_COMP_lpi_1_dfm_4);
      COMP_i_0_1_lpi_1_dfm_6 <= COMP_i_0_1_lpi_1_dfm_5;
      pe_x_reg_0_lpi_1_dfm_4 <= pe_x_reg_0_lpi_1_dfm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exit_for_for_for_1_lpi_1_dfm_1_st_4 <= 1'b0;
    end
    else if ( core_wen & (~(lfst_exit_for_for_for_1_lpi_1_dfm_st_1_0 & lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1))
        & main_stage_0_2 ) begin
      exit_for_for_for_1_lpi_1_dfm_1_st_4 <= MUX_s_1_2_2(exitL_exit_COL_1_COMP_lpi_1_dfm_4,
          exit_for_for_for_1_lpi_1_dfm_1_st_3, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pe_y_reg_value_15_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_14_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_13_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_12_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_11_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_10_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_9_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_8_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_7_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_6_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_5_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_4_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_3_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_2_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_1_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_0_63_32_lpi_2 <= 32'b0;
      pe_y_reg_value_15_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_14_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_13_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_12_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_11_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_10_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_9_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_8_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_7_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_6_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_5_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_4_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_3_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_2_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_1_31_0_lpi_2 <= 32'b0;
      pe_y_reg_value_0_31_0_lpi_2 <= 32'b0;
    end
    else if ( pe_y_reg_value_and_cse ) begin
      pe_y_reg_value_15_63_32_lpi_2 <= pe_y_reg_value_15_63_32_sva_1_mx0;
      pe_y_reg_value_14_63_32_lpi_2 <= pe_y_reg_value_14_63_32_sva_1_mx0;
      pe_y_reg_value_13_63_32_lpi_2 <= pe_y_reg_value_13_63_32_sva_1_mx0;
      pe_y_reg_value_12_63_32_lpi_2 <= pe_y_reg_value_12_63_32_sva_1_mx0;
      pe_y_reg_value_11_63_32_lpi_2 <= pe_y_reg_value_11_63_32_sva_1_mx0;
      pe_y_reg_value_10_63_32_lpi_2 <= pe_y_reg_value_10_63_32_sva_1_mx0;
      pe_y_reg_value_9_63_32_lpi_2 <= pe_y_reg_value_9_63_32_sva_1_mx0;
      pe_y_reg_value_8_63_32_lpi_2 <= pe_y_reg_value_8_63_32_sva_1_mx0;
      pe_y_reg_value_7_63_32_lpi_2 <= pe_y_reg_value_7_63_32_sva_1_mx0;
      pe_y_reg_value_6_63_32_lpi_2 <= pe_y_reg_value_6_63_32_sva_1_mx0;
      pe_y_reg_value_5_63_32_lpi_2 <= pe_y_reg_value_5_63_32_sva_1_mx0;
      pe_y_reg_value_4_63_32_lpi_2 <= pe_y_reg_value_4_63_32_sva_1_mx0;
      pe_y_reg_value_3_63_32_lpi_2 <= pe_y_reg_value_3_63_32_sva_1_mx0;
      pe_y_reg_value_2_63_32_lpi_2 <= pe_y_reg_value_2_63_32_sva_1_mx0;
      pe_y_reg_value_1_63_32_lpi_2 <= pe_y_reg_value_1_63_32_sva_1_mx0;
      pe_y_reg_value_0_63_32_lpi_2 <= pe_y_reg_value_0_63_32_sva_1_mx0;
      pe_y_reg_value_15_31_0_lpi_2 <= pe_y_reg_value_15_31_0_sva_1_mx0;
      pe_y_reg_value_14_31_0_lpi_2 <= pe_y_reg_value_14_31_0_sva_1_mx0;
      pe_y_reg_value_13_31_0_lpi_2 <= pe_y_reg_value_13_31_0_sva_1_mx0;
      pe_y_reg_value_12_31_0_lpi_2 <= pe_y_reg_value_12_31_0_sva_1_mx0;
      pe_y_reg_value_11_31_0_lpi_2 <= pe_y_reg_value_11_31_0_sva_1_mx0;
      pe_y_reg_value_10_31_0_lpi_2 <= pe_y_reg_value_10_31_0_sva_1_mx0;
      pe_y_reg_value_9_31_0_lpi_2 <= pe_y_reg_value_9_31_0_sva_1_mx0;
      pe_y_reg_value_8_31_0_lpi_2 <= pe_y_reg_value_8_31_0_sva_1_mx0;
      pe_y_reg_value_7_31_0_lpi_2 <= pe_y_reg_value_7_31_0_sva_1_mx0;
      pe_y_reg_value_6_31_0_lpi_2 <= pe_y_reg_value_6_31_0_sva_1_mx0;
      pe_y_reg_value_5_31_0_lpi_2 <= pe_y_reg_value_5_31_0_sva_1_mx0;
      pe_y_reg_value_4_31_0_lpi_2 <= pe_y_reg_value_4_31_0_sva_1_mx0;
      pe_y_reg_value_3_31_0_lpi_2 <= pe_y_reg_value_3_31_0_sva_1_mx0;
      pe_y_reg_value_2_31_0_lpi_2 <= pe_y_reg_value_2_31_0_sva_1_mx0;
      pe_y_reg_value_1_31_0_lpi_2 <= pe_y_reg_value_1_31_0_sva_1_mx0;
      pe_y_reg_value_0_31_0_lpi_2 <= pe_y_reg_value_0_31_0_sva_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_lo_conc_1_itm_2_5_1 <= 1'b0;
      reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp <= 1'b0;
      reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp_1 <= 3'b0;
    end
    else if ( PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_and_cse ) begin
      PackedStencil_DTYPE_2U_1U_1U_1U_operator_4_lo_conc_1_itm_2_5_1 <= out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1;
      reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp <= reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_itm;
      reg_for_for_for_1_k_slc_for_for_for_1_k_4_0_3_0_ssc_2_tmp_1 <= reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_1_itm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 <= 1'b0;
      lfst_exit_for_for_for_1_lpi_1_dfm_st_2_0_1 <= 1'b0;
      for_for_for_1_equal_tmp_10 <= 1'b0;
      for_for_for_1_equal_tmp_12 <= 1'b0;
      lfst_exit_for_for_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( for_for_for_1_and_291_cse ) begin
      lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 <= lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1;
      lfst_exit_for_for_for_1_lpi_1_dfm_st_2_0_1 <= lfst_exit_for_for_for_1_lpi_1_dfm_st_1_0;
      for_for_for_1_equal_tmp_10 <= for_for_for_1_equal_tmp_2;
      for_for_for_1_equal_tmp_12 <= for_for_for_1_equal_tmp_5;
      lfst_exit_for_for_1_lpi_1_dfm_4 <= lfst_exit_for_for_1_lpi_1_dfm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_row_slc_for_for_row_6_0_5_0_1_itm_3 <= 6'b0;
      WX_if_1_acc_decb_sva_1_3_1_1 <= 3'b0;
    end
    else if ( for_for_row_and_cse ) begin
      for_for_row_slc_for_for_row_6_0_5_0_1_itm_3 <= for_for_row_6_0_lpi_1_dfm[5:0];
      WX_if_1_acc_decb_sva_1_3_1_1 <= MUX_v_3_2_2(WX_if_1_acc_decb_sva_3_1_mx0w0,
          WX_if_1_acc_decb_sva_3_1, and_233_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exit_WY_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_65 | or_dcpl_38)) ) begin
      exit_WY_sva_2 <= ~ WY_acc_tmp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_i_0_15_lpi_1 <= 1'b0;
      COMP_i_0_14_lpi_1 <= 1'b0;
      COMP_i_0_13_lpi_1 <= 1'b0;
      COMP_i_0_12_lpi_1 <= 1'b0;
      COMP_i_0_11_lpi_1 <= 1'b0;
      COMP_i_0_10_lpi_1 <= 1'b0;
      COMP_i_0_9_lpi_1 <= 1'b0;
      COMP_i_0_8_lpi_1 <= 1'b0;
      COMP_i_0_7_lpi_1 <= 1'b0;
      COMP_i_0_6_lpi_1 <= 1'b0;
      COMP_i_0_5_lpi_1 <= 1'b0;
      COMP_i_0_4_lpi_1 <= 1'b0;
      COMP_i_0_3_lpi_1 <= 1'b0;
      COMP_i_0_2_lpi_1 <= 1'b0;
      COMP_i_0_1_lpi_1 <= 1'b0;
      COMP_i_0_lpi_1 <= 1'b0;
      exitL_exit_COL_1_COMP_lpi_1 <= 1'b0;
      lfst_exit_WX_1_lpi_1 <= 1'b0;
      exitL_exit_COL_1_COMP_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( COMP_i_and_cse ) begin
      COMP_i_0_15_lpi_1 <= ~ COMP_i_0_15_lpi_1_dfm;
      COMP_i_0_14_lpi_1 <= ~ COMP_i_0_14_lpi_1_dfm;
      COMP_i_0_13_lpi_1 <= ~ COMP_i_0_13_lpi_1_dfm;
      COMP_i_0_12_lpi_1 <= ~ COMP_i_0_12_lpi_1_dfm;
      COMP_i_0_11_lpi_1 <= ~ COMP_i_0_11_lpi_1_dfm;
      COMP_i_0_10_lpi_1 <= ~ COMP_i_0_10_lpi_1_dfm;
      COMP_i_0_9_lpi_1 <= ~ COMP_i_0_9_lpi_1_dfm;
      COMP_i_0_8_lpi_1 <= ~ COMP_i_0_8_lpi_1_dfm;
      COMP_i_0_7_lpi_1 <= ~ COMP_i_0_7_lpi_1_dfm;
      COMP_i_0_6_lpi_1 <= ~ COMP_i_0_6_lpi_1_dfm;
      COMP_i_0_5_lpi_1 <= ~ COMP_i_0_5_lpi_1_dfm;
      COMP_i_0_4_lpi_1 <= ~ COMP_i_0_4_lpi_1_dfm;
      COMP_i_0_3_lpi_1 <= ~ COMP_i_0_3_lpi_1_dfm;
      COMP_i_0_2_lpi_1 <= ~ COMP_i_0_2_lpi_1_dfm;
      COMP_i_0_1_lpi_1 <= ~ COMP_i_0_1_lpi_1_dfm;
      COMP_i_0_lpi_1 <= ~ COMP_i_0_lpi_1_dfm;
      exitL_exit_COL_1_COMP_lpi_1 <= COMP_and_13_tmp;
      lfst_exit_WX_1_lpi_1 <= ~ exit_WX_lpi_1_dfm_1;
      exitL_exit_COL_1_COMP_lpi_1_dfm_4 <= exitL_exit_COL_1_COMP_lpi_1_dfm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      WX_wx_1_0_lpi_3 <= 2'b0;
    end
    else if ( (WY_mux_6_tmp==2'b01) & core_wen & or_71_cse ) begin
      WX_wx_1_0_lpi_3 <= for_for_for_1_for_for_for_1_for_for_for_1_mux1h_1_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_1_k_4_0_lpi_1_3_0_1 <= 4'b0;
    end
    else if ( (mux_201_nl) & core_wen ) begin
      for_for_for_1_k_4_0_lpi_1_3_0_1 <= MUX_v_4_2_2((WY_WY_and_2_nl), (for_for_for_1_acc_1_tmp[3:0]),
          for_for_for_1_and_97_cse);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_1_for_q_0_lpi_2 <= 1'b0;
    end
    else if ( core_wen & (for_for_for_1_nor_dfs | for_for_for_1_and_97_cse | for_for_for_1_asn_rgt_4)
        ) begin
      for_for_for_1_for_q_0_lpi_2 <= MUX1HOT_s_1_3_2((WY_WY_and_3_nl), (and_55_nl),
          (~ for_for_for_1_for_q_0_lpi_2), {for_for_for_1_nor_dfs , for_for_for_1_and_97_cse
          , for_for_for_1_asn_rgt_4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      WY_wy_1_0_lpi_3 <= 2'b0;
      for_for_for_1_nor_dfs_5 <= 1'b0;
      unequal_tmp_5 <= 1'b0;
    end
    else if ( WY_wy_and_cse ) begin
      WY_wy_1_0_lpi_3 <= MUX_v_2_2_2(2'b00, (mux_203_nl), (nor_64_nl));
      for_for_for_1_nor_dfs_5 <= for_for_for_1_nor_dfs;
      unequal_tmp_5 <= unequal_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_row_6_0_lpi_3 <= 7'b0;
      for_ko_2_0_lpi_1_1_0_1 <= 2'b0;
    end
    else if ( for_for_row_and_1_cse ) begin
      for_for_row_6_0_lpi_3 <= MUX1HOT_v_7_3_2(for_for_row_6_0_lpi_1_dfm, (signext_7_1(for_acc_2_tmp[2])),
          for_for_acc_1_tmp, {(for_for_for_1_nand_nl) , (for_for_for_1_and_nl) ,
          (for_for_for_1_and_166_nl)});
      for_ko_2_0_lpi_1_1_0_1 <= MUX_v_2_2_2(for_ko_2_0_lpi_1_dfm_1_0, (for_acc_2_tmp[1:0]),
          and_232_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out_tmp_value_0_31_0_lpi_2 <= 32'b0;
    end
    else if ( (~ (mux_206_nl)) & core_wen ) begin
      out_tmp_value_0_31_0_lpi_2 <= MUX_v_32_2_2(out_tmp_value_0_31_0_lpi_1_mx0w0,
          (and_59_nl), main_stage_0_3);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_33_itm_2 <= 32'b0;
    end
    else if ( (mux_208_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_33_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_15_31_0_sva_1_mx0, out_tmp_value_15_31_0_lpi_1_dfm_mx0w0,
          ({{16{COL_7_COMP_tmp_acc_psp_sva[15]}}, COL_7_COMP_tmp_acc_psp_sva}), pe_y_reg_value_6_63_32_lpi_1_dfm_mx0,
          {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6) , and_dcpl_70 , and_dcpl_71});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_row_6_0_lpi_1_dfm_7_6_1 <= 1'b0;
    end
    else if ( core_wen & or_395_cse & for_for_for_1_nor_dfs_6 & (~ lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1)
        & (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5==2'b00) & (~ unequal_tmp_6) &
        main_stage_0_3 ) begin
      for_for_row_6_0_lpi_1_dfm_7_6_1 <= for_for_row_6_0_lpi_1_dfm_6_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_32_itm_2 <= 32'b0;
    end
    else if ( (mux_210_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_32_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_15_63_32_sva_1_mx0, out_tmp_value_15_63_32_lpi_1_dfm_mx0w0,
          pe_y_reg_value_6_31_0_lpi_1_dfm_mx0, ({{16{COL_7_COMP_tmp_acc_psp_sva[15]}},
          COL_7_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_70 , and_dcpl_71});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_31_itm_2 <= 32'b0;
    end
    else if ( (mux_212_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_31_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_14_31_0_sva_1_mx0, out_tmp_value_14_31_0_lpi_1_dfm_mx0w0,
          ({{16{COL_6_COMP_tmp_acc_psp_sva[15]}}, COL_6_COMP_tmp_acc_psp_sva}), pe_y_reg_value_5_63_32_lpi_1_dfm_mx0,
          {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6) , and_dcpl_72 , and_dcpl_73});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_30_itm_2 <= 32'b0;
    end
    else if ( (mux_214_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_30_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_14_63_32_sva_1_mx0, out_tmp_value_14_63_32_lpi_1_dfm_mx0w0,
          pe_y_reg_value_5_31_0_lpi_1_dfm_mx0, ({{16{COL_6_COMP_tmp_acc_psp_sva[15]}},
          COL_6_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_72 , and_dcpl_73});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_29_itm_2 <= 32'b0;
    end
    else if ( (mux_216_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_29_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_13_31_0_sva_1_mx0, out_tmp_value_13_31_0_lpi_1_dfm_mx0w0,
          pe_y_reg_value_4_31_0_lpi_1_dfm_mx0, ({{16{COL_5_COMP_tmp_acc_psp_sva[15]}},
          COL_5_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_74 , and_dcpl_75});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_28_itm_2 <= 32'b0;
    end
    else if ( (mux_218_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_28_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_13_63_32_sva_1_mx0, out_tmp_value_13_63_32_lpi_1_dfm_mx0w0,
          ({{16{COL_4_COMP_tmp_acc_psp_sva[15]}}, COL_4_COMP_tmp_acc_psp_sva}), pe_y_reg_value_3_63_32_lpi_1_dfm_mx0,
          {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6) , and_dcpl_76 , and_dcpl_77});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_27_itm_2 <= 32'b0;
    end
    else if ( (mux_220_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_27_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_12_31_0_sva_1_mx0, out_tmp_value_12_31_0_lpi_1_dfm_mx0w0,
          pe_y_reg_value_3_31_0_lpi_1_dfm_mx0, ({{16{COL_4_COMP_tmp_acc_psp_sva[15]}},
          COL_4_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_76 , and_dcpl_77});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_26_itm_2 <= 32'b0;
    end
    else if ( (mux_222_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_26_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_12_63_32_sva_1_mx0, out_tmp_value_12_63_32_lpi_1_dfm_mx0w0,
          ({{16{COL_3_COMP_tmp_acc_psp_sva[15]}}, COL_3_COMP_tmp_acc_psp_sva}), pe_y_reg_value_2_63_32_lpi_1_dfm_mx0,
          {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6) , and_dcpl_78 , and_dcpl_79});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_25_itm_2 <= 32'b0;
    end
    else if ( (mux_224_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_25_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_11_31_0_sva_1_mx0, out_tmp_value_11_31_0_lpi_1_dfm_mx0w0,
          pe_y_reg_value_2_31_0_lpi_1_dfm_mx0, ({{16{COL_3_COMP_tmp_acc_psp_sva[15]}},
          COL_3_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_78 , and_dcpl_79});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_24_itm_2 <= 32'b0;
    end
    else if ( (mux_226_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_24_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_11_63_32_sva_1_mx0, out_tmp_value_11_63_32_lpi_1_dfm_mx0w0,
          ({{16{COL_16_COMP_tmp_acc_psp_sva[15]}}, COL_16_COMP_tmp_acc_psp_sva}),
          pe_y_reg_value_15_63_32_lpi_1_dfm_mx0, {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_80 , and_dcpl_81});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_23_itm_2 <= 32'b0;
    end
    else if ( (mux_228_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_23_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_10_31_0_sva_1_mx0, out_tmp_value_10_31_0_lpi_1_dfm_mx0w0,
          pe_y_reg_value_15_31_0_lpi_1_dfm_mx0, ({{16{COL_16_COMP_tmp_acc_psp_sva[15]}},
          COL_16_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_80 , and_dcpl_81});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_22_itm_2 <= 32'b0;
    end
    else if ( (mux_230_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_22_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_10_63_32_sva_1_mx0, out_tmp_value_10_63_32_lpi_1_dfm_mx0w0,
          ({{16{COL_15_COMP_tmp_acc_psp_sva[15]}}, COL_15_COMP_tmp_acc_psp_sva}),
          pe_y_reg_value_14_63_32_lpi_1_dfm_mx0, {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_82 , and_dcpl_83});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_21_itm_2 <= 32'b0;
    end
    else if ( (mux_232_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_21_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_9_31_0_sva_1_mx0, out_tmp_value_9_31_0_lpi_1_dfm,
          pe_y_reg_value_14_31_0_lpi_1_dfm_mx0, ({{16{COL_15_COMP_tmp_acc_psp_sva[15]}},
          COL_15_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_82 , and_dcpl_83});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_20_itm_2 <= 32'b0;
    end
    else if ( (mux_234_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_20_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_9_63_32_sva_1_mx0, out_tmp_value_9_63_32_lpi_1_dfm,
          ({{16{COL_14_COMP_tmp_acc_psp_sva[15]}}, COL_14_COMP_tmp_acc_psp_sva}),
          pe_y_reg_value_13_63_32_lpi_1_dfm_mx0, {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_84 , and_dcpl_85});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_19_itm_2 <= 32'b0;
    end
    else if ( (mux_236_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_19_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_8_31_0_sva_1_mx0, out_tmp_value_8_31_0_lpi_1_dfm,
          ({{16{COL_13_COMP_tmp_acc_psp_sva[15]}}, COL_13_COMP_tmp_acc_psp_sva}),
          pe_y_reg_value_12_63_32_lpi_1_dfm_mx0, {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_86 , and_dcpl_87});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_18_itm_2 <= 32'b0;
    end
    else if ( (mux_238_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_18_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_8_63_32_sva_1_mx0, out_tmp_value_8_63_32_lpi_1_dfm,
          pe_y_reg_value_12_31_0_lpi_1_dfm_mx0, ({{16{COL_13_COMP_tmp_acc_psp_sva[15]}},
          COL_13_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_86 , and_dcpl_87});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_17_itm_2 <= 32'b0;
    end
    else if ( (mux_240_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_17_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_7_31_0_sva_1_mx0, out_tmp_value_7_31_0_lpi_1_dfm,
          ({{16{COL_12_COMP_tmp_acc_psp_sva[15]}}, COL_12_COMP_tmp_acc_psp_sva}),
          pe_y_reg_value_11_63_32_lpi_1_dfm_mx0, {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_88 , and_dcpl_89});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_16_itm_2 <= 32'b0;
    end
    else if ( (mux_242_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_16_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_7_63_32_sva_1_mx0, out_tmp_value_7_63_32_lpi_1_dfm,
          pe_y_reg_value_11_31_0_lpi_1_dfm_mx0, ({{16{COL_12_COMP_tmp_acc_psp_sva[15]}},
          COL_12_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_88 , and_dcpl_89});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_15_itm_2 <= 32'b0;
    end
    else if ( (mux_244_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_15_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_6_31_0_sva_1_mx0, out_tmp_value_6_31_0_lpi_1_dfm,
          ({{16{COL_11_COMP_tmp_acc_psp_sva[15]}}, COL_11_COMP_tmp_acc_psp_sva}),
          pe_y_reg_value_10_63_32_lpi_1_dfm_mx0, {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_90 , and_dcpl_91});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_14_itm_2 <= 32'b0;
    end
    else if ( (mux_246_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_14_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_6_63_32_sva_1_mx0, out_tmp_value_6_63_32_lpi_1_dfm,
          pe_y_reg_value_10_31_0_lpi_1_dfm_mx0, ({{16{COL_11_COMP_tmp_acc_psp_sva[15]}},
          COL_11_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_90 , and_dcpl_91});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_13_itm_2 <= 32'b0;
    end
    else if ( (mux_248_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_13_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_5_31_0_sva_1_mx0, out_tmp_value_5_31_0_lpi_1_dfm,
          ({{16{COL_2_COMP_tmp_acc_psp_sva[15]}}, COL_2_COMP_tmp_acc_psp_sva}), pe_y_reg_value_1_63_32_lpi_1_dfm_mx0,
          {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6) , and_dcpl_92 , and_dcpl_93});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_12_itm_2 <= 32'b0;
    end
    else if ( (mux_250_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_12_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_5_63_32_sva_1_mx0, out_tmp_value_5_63_32_lpi_1_dfm,
          pe_y_reg_value_1_31_0_lpi_1_dfm_mx0, ({{16{COL_2_COMP_tmp_acc_psp_sva[15]}},
          COL_2_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_92 , and_dcpl_93});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_11_itm_2 <= 32'b0;
    end
    else if ( (mux_252_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_11_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_4_31_0_sva_1_mx0, out_tmp_value_4_31_0_lpi_1_dfm,
          ({{16{COL_1_COMP_tmp_acc_psp_sva[15]}}, COL_1_COMP_tmp_acc_psp_sva}), pe_y_reg_value_0_63_32_lpi_1_dfm_mx0,
          {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6) , and_dcpl_94 , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_10_itm_2 <= 32'b0;
    end
    else if ( (mux_254_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_10_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_4_63_32_sva_1_mx0, out_tmp_value_4_63_32_lpi_1_dfm,
          pe_y_reg_value_0_31_0_lpi_1_dfm_mx0, ({{16{COL_1_COMP_tmp_acc_psp_sva[15]}},
          COL_1_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_94 , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_9_itm_2 <= 32'b0;
    end
    else if ( (mux_256_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_9_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_3_31_0_sva_1_mx0, out_tmp_value_3_31_0_lpi_1_dfm,
          ({{16{COL_10_COMP_tmp_acc_psp_sva[15]}}, COL_10_COMP_tmp_acc_psp_sva}),
          pe_y_reg_value_9_63_32_lpi_1_dfm_mx0, {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_96 , and_dcpl_97});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_8_itm_2 <= 32'b0;
    end
    else if ( (mux_258_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_8_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_3_63_32_sva_1_mx0, out_tmp_value_3_63_32_lpi_1_dfm,
          pe_y_reg_value_9_31_0_lpi_1_dfm_mx0, ({{16{COL_10_COMP_tmp_acc_psp_sva[15]}},
          COL_10_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_96 , and_dcpl_97});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_7_itm_2 <= 32'b0;
    end
    else if ( (mux_260_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_7_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_2_31_0_sva_1_mx0, out_tmp_value_2_31_0_lpi_1_dfm,
          ({{16{COL_9_COMP_tmp_acc_psp_sva[15]}}, COL_9_COMP_tmp_acc_psp_sva}), pe_y_reg_value_8_63_32_lpi_1_dfm_mx0,
          {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6) , and_dcpl_98 , and_dcpl_99});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_6_itm_2 <= 32'b0;
    end
    else if ( (mux_262_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_6_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_2_63_32_sva_1_mx0, out_tmp_value_2_63_32_lpi_1_dfm,
          pe_y_reg_value_8_31_0_lpi_1_dfm_mx0, ({{16{COL_9_COMP_tmp_acc_psp_sva[15]}},
          COL_9_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_98 , and_dcpl_99});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_5_itm_2 <= 32'b0;
    end
    else if ( (mux_264_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_5_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_1_31_0_sva_1_mx0, out_tmp_value_1_31_0_lpi_1_dfm_mx0w0,
          ({{16{COL_8_COMP_tmp_acc_psp_sva[15]}}, COL_8_COMP_tmp_acc_psp_sva}), pe_y_reg_value_7_63_32_lpi_1_dfm_mx0,
          {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6) , and_dcpl_100 , and_dcpl_101});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_4_itm_2 <= 32'b0;
    end
    else if ( (mux_266_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_4_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_1_63_32_sva_1_mx0, out_tmp_value_1_63_32_lpi_1_dfm_mx0w0,
          pe_y_reg_value_7_31_0_lpi_1_dfm_mx0, ({{16{COL_8_COMP_tmp_acc_psp_sva[15]}},
          COL_8_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_100 , and_dcpl_101});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_3_itm_2 <= 32'b0;
    end
    else if ( (mux_268_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_3_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_0_31_0_sva_1_mx0, out_tmp_value_0_31_0_lpi_1_dfm_mx0w0,
          ({{16{COL_5_COMP_tmp_acc_psp_sva[15]}}, COL_5_COMP_tmp_acc_psp_sva}), pe_y_reg_value_4_63_32_lpi_1_dfm_mx0,
          {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6) , and_dcpl_74 , and_dcpl_75});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_mux_2_itm_2 <= 32'b0;
    end
    else if ( (mux_270_nl) & core_wen & and_dcpl_15 ) begin
      COMP_mux_2_itm_2 <= MUX1HOT_v_32_4_2(pe_y_reg_value_0_63_32_sva_1_mx0, out_tmp_value_0_63_32_lpi_1_dfm_mx0w0,
          pe_y_reg_value_13_31_0_lpi_1_dfm_mx0, ({{16{COL_14_COMP_tmp_acc_psp_sva[15]}},
          COL_14_COMP_tmp_acc_psp_sva}), {and_dcpl_68 , (~ COMP_and_13_mdf_sva_6)
          , and_dcpl_84 , and_dcpl_85});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out_tmp_value_15_31_0_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_15_63_32_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_14_31_0_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_14_63_32_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_13_31_0_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_13_63_32_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_12_31_0_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_12_63_32_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_11_31_0_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_11_63_32_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_10_31_0_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_10_63_32_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_1_31_0_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_1_63_32_lpi_1_dfm_11 <= 32'b0;
      out_tmp_value_0_31_0_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_0_63_32_lpi_1_dfm_11 <= 32'b0;
    end
    else if ( out_tmp_value_and_1_cse ) begin
      out_tmp_value_15_31_0_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_15_31_0_lpi_1_dfm_mx0w0,
          out_tmp_value_8_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_15_63_32_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_15_63_32_lpi_1_dfm_mx0w0,
          out_tmp_value_9_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_14_31_0_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_14_31_0_lpi_1_dfm_mx0w0,
          out_tmp_value_6_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_14_63_32_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_14_63_32_lpi_1_dfm_mx0w0,
          out_tmp_value_7_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_13_31_0_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_13_31_0_lpi_1_dfm_mx0w0,
          out_tmp_value_4_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_13_63_32_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_13_63_32_lpi_1_dfm_mx0w0,
          out_tmp_value_5_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_12_31_0_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_12_31_0_lpi_1_dfm_mx0w0,
          out_tmp_value_2_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_12_63_32_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_12_63_32_lpi_1_dfm_mx0w0,
          out_tmp_value_3_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_11_31_0_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_11_31_0_lpi_1_dfm_mx0w0,
          out_tmp_value_14_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_11_63_32_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_11_63_32_lpi_1_dfm_mx0w0,
          out_tmp_value_15_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_10_31_0_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_10_31_0_lpi_1_dfm_mx0w0,
          out_tmp_value_12_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_10_63_32_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_10_63_32_lpi_1_dfm_mx0w0,
          out_tmp_value_13_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_1_31_0_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_1_31_0_lpi_1_dfm_mx0w0,
          out_tmp_value_10_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_1_63_32_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_1_63_32_lpi_1_dfm_mx0w0,
          out_tmp_value_11_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_0_31_0_lpi_1_dfm_10 <= MUX_v_32_2_2(out_tmp_value_0_31_0_lpi_1_dfm_mx0w0,
          out_tmp_value_0_63_32_lpi_1_mx0w0, and_dcpl_66);
      out_tmp_value_0_63_32_lpi_1_dfm_11 <= MUX_v_32_2_2(out_tmp_value_0_63_32_lpi_1_dfm_mx0w0,
          out_tmp_value_1_63_32_lpi_1_mx0w0, and_dcpl_66);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out_tmp_value_15_31_0_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_15_63_32_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_14_31_0_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_14_63_32_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_13_31_0_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_13_63_32_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_12_31_0_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_12_63_32_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_11_31_0_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_11_63_32_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_10_31_0_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_10_63_32_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_1_31_0_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_1_63_32_lpi_1_dfm_10 <= 32'b0;
      out_tmp_value_0_63_32_lpi_1_dfm_10 <= 32'b0;
    end
    else if ( out_tmp_value_and_2_cse ) begin
      out_tmp_value_15_31_0_lpi_1_dfm_10 <= MUX_v_32_2_2((and_89_nl), out_tmp_value_8_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_15_63_32_lpi_1_dfm_10 <= MUX_v_32_2_2((and_88_nl), out_tmp_value_9_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_14_31_0_lpi_1_dfm_10 <= MUX_v_32_2_2((and_87_nl), out_tmp_value_6_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_14_63_32_lpi_1_dfm_10 <= MUX_v_32_2_2((and_86_nl), out_tmp_value_7_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_13_31_0_lpi_1_dfm_10 <= MUX_v_32_2_2((and_85_nl), out_tmp_value_4_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_13_63_32_lpi_1_dfm_10 <= MUX_v_32_2_2((and_84_nl), out_tmp_value_5_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_12_31_0_lpi_1_dfm_10 <= MUX_v_32_2_2((and_83_nl), out_tmp_value_2_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_12_63_32_lpi_1_dfm_10 <= MUX_v_32_2_2((and_82_nl), out_tmp_value_3_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_11_31_0_lpi_1_dfm_10 <= MUX_v_32_2_2((and_81_nl), out_tmp_value_14_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_11_63_32_lpi_1_dfm_10 <= MUX_v_32_2_2((and_80_nl), out_tmp_value_15_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_10_31_0_lpi_1_dfm_10 <= MUX_v_32_2_2((and_79_nl), out_tmp_value_12_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_10_63_32_lpi_1_dfm_10 <= MUX_v_32_2_2((and_78_nl), out_tmp_value_13_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_1_31_0_lpi_1_dfm_10 <= MUX_v_32_2_2((and_61_nl), out_tmp_value_10_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_1_63_32_lpi_1_dfm_10 <= MUX_v_32_2_2((and_60_nl), out_tmp_value_11_31_0_lpi_1_mx0w0,
          and_dcpl_66);
      out_tmp_value_0_63_32_lpi_1_dfm_10 <= MUX_v_32_2_2((and_58_nl), out_tmp_value_1_31_0_lpi_1_mx0w0,
          and_dcpl_66);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out_tmp_value_9_31_0_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_9_63_32_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_8_31_0_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_8_63_32_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_7_31_0_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_7_63_32_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_6_31_0_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_6_63_32_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_5_31_0_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_5_63_32_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_4_31_0_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_4_63_32_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_3_31_0_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_3_63_32_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_2_31_0_lpi_1_dfm_13 <= 32'b0;
      out_tmp_value_2_63_32_lpi_1_dfm_13 <= 32'b0;
    end
    else if ( out_tmp_value_and_25_cse ) begin
      out_tmp_value_9_31_0_lpi_1_dfm_13 <= out_tmp_value_9_31_0_lpi_1_dfm;
      out_tmp_value_9_63_32_lpi_1_dfm_13 <= out_tmp_value_9_63_32_lpi_1_dfm;
      out_tmp_value_8_31_0_lpi_1_dfm_13 <= out_tmp_value_8_31_0_lpi_1_dfm;
      out_tmp_value_8_63_32_lpi_1_dfm_13 <= out_tmp_value_8_63_32_lpi_1_dfm;
      out_tmp_value_7_31_0_lpi_1_dfm_13 <= out_tmp_value_7_31_0_lpi_1_dfm;
      out_tmp_value_7_63_32_lpi_1_dfm_13 <= out_tmp_value_7_63_32_lpi_1_dfm;
      out_tmp_value_6_31_0_lpi_1_dfm_13 <= out_tmp_value_6_31_0_lpi_1_dfm;
      out_tmp_value_6_63_32_lpi_1_dfm_13 <= out_tmp_value_6_63_32_lpi_1_dfm;
      out_tmp_value_5_31_0_lpi_1_dfm_13 <= out_tmp_value_5_31_0_lpi_1_dfm;
      out_tmp_value_5_63_32_lpi_1_dfm_13 <= out_tmp_value_5_63_32_lpi_1_dfm;
      out_tmp_value_4_31_0_lpi_1_dfm_13 <= out_tmp_value_4_31_0_lpi_1_dfm;
      out_tmp_value_4_63_32_lpi_1_dfm_13 <= out_tmp_value_4_63_32_lpi_1_dfm;
      out_tmp_value_3_31_0_lpi_1_dfm_13 <= out_tmp_value_3_31_0_lpi_1_dfm;
      out_tmp_value_3_63_32_lpi_1_dfm_13 <= out_tmp_value_3_63_32_lpi_1_dfm;
      out_tmp_value_2_31_0_lpi_1_dfm_13 <= out_tmp_value_2_31_0_lpi_1_dfm;
      out_tmp_value_2_63_32_lpi_1_dfm_13 <= out_tmp_value_2_63_32_lpi_1_dfm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out_tmp_value_9_31_0_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_9_63_32_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_8_31_0_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_8_63_32_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_7_31_0_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_7_63_32_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_6_31_0_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_6_63_32_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_5_31_0_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_5_63_32_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_4_31_0_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_4_63_32_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_3_31_0_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_3_63_32_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_2_31_0_lpi_1_dfm_12 <= 32'b0;
      out_tmp_value_2_63_32_lpi_1_dfm_12 <= 32'b0;
    end
    else if ( out_tmp_value_and_26_cse ) begin
      out_tmp_value_9_31_0_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_9_31_0_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_9_63_32_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_9_63_32_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_8_31_0_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_8_31_0_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_8_63_32_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_8_63_32_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_7_31_0_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_7_31_0_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_7_63_32_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_7_63_32_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_6_31_0_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_6_31_0_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_6_63_32_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_6_63_32_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_5_31_0_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_5_31_0_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_5_63_32_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_5_63_32_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_4_31_0_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_4_31_0_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_4_63_32_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_4_63_32_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_3_31_0_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_3_31_0_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_3_63_32_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_3_63_32_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_2_31_0_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_2_31_0_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
      out_tmp_value_2_63_32_lpi_1_dfm_12 <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          out_tmp_value_2_63_32_lpi_1_dfm, for_for_row_6_0_lpi_1_dfm_6_6_1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exit_for_for_for_1_lpi_1_dfm_10_1_1 <= 1'b0;
      COMP_and_13_mdf_sva_7 <= 1'b0;
      for_for_for_1_equal_tmp_13 <= 1'b0;
      unequal_tmp_7 <= 1'b0;
      for_for_for_1_nor_dfs_7 <= 1'b0;
    end
    else if ( for_for_for_1_and_293_cse ) begin
      lfst_exit_for_for_for_1_lpi_1_dfm_10_1_1 <= lfst_exit_for_for_for_1_lpi_1_dfm_9_1_1;
      COMP_and_13_mdf_sva_7 <= COMP_and_13_mdf_sva_6;
      for_for_for_1_equal_tmp_13 <= for_for_for_1_equal_tmp_12;
      unequal_tmp_7 <= unequal_tmp_6;
      for_for_for_1_nor_dfs_7 <= for_for_for_1_nor_dfs_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000
          <= 16'b0;
    end
    else if ( (~((out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1
        | (reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_1_itm[1:0]!=2'b00))
        & (reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_1_itm[2])))
        & (~ lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1) & main_stage_0_2 & core_wen
        ) begin
      COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_COL_1_PackedStencil_DTYPE_2U_1U_1U_1U_operator_1_slc_weight_buf_value_64_63_0_cse_47_0_COL_1_PackedStencil000000
          <= MUX_v_16_9_2((mux1h_45_nl), (mux1h_44_nl), (mux1h_43_nl), (mux1h_42_nl),
          (mux1h_41_nl), (mux1h_40_nl), (mux1h_39_nl), (mux1h_38_nl), (mux1h_nl),
          {reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_1_itm
          , out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exit_for_for_for_1_lpi_1_dfm_1_st_3 <= 1'b0;
    end
    else if ( core_wen & and_dcpl_27 ) begin
      exit_for_for_for_1_lpi_1_dfm_1_st_3 <= exit_for_for_for_1_lpi_1_dfm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exit_for_for_for_1_lpi_1_dfm_1_st_4 <= 2'b0;
      WX_unequal_tmp_5 <= 1'b0;
      COMP_i_0_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_2_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_3_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_4_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_5_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_6_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_7_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_8_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_9_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_10_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_11_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_12_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_13_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_14_lpi_1_dfm_5 <= 1'b0;
      COMP_i_0_15_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( for_for_for_1_and_299_cse ) begin
      lfst_exit_for_for_for_1_lpi_1_dfm_1_st_4 <= WY_mux_3_cse;
      WX_unequal_tmp_5 <= (WX_wx_1_0_lpi_1_dfm!=2'b00);
      COMP_i_0_lpi_1_dfm_5 <= COMP_i_0_lpi_1_dfm;
      COMP_i_0_2_lpi_1_dfm_5 <= COMP_i_0_2_lpi_1_dfm;
      COMP_i_0_3_lpi_1_dfm_5 <= COMP_i_0_3_lpi_1_dfm;
      COMP_i_0_4_lpi_1_dfm_5 <= COMP_i_0_4_lpi_1_dfm;
      COMP_i_0_5_lpi_1_dfm_5 <= COMP_i_0_5_lpi_1_dfm;
      COMP_i_0_6_lpi_1_dfm_5 <= COMP_i_0_6_lpi_1_dfm;
      COMP_i_0_7_lpi_1_dfm_5 <= COMP_i_0_7_lpi_1_dfm;
      COMP_i_0_8_lpi_1_dfm_5 <= COMP_i_0_8_lpi_1_dfm;
      COMP_i_0_9_lpi_1_dfm_5 <= COMP_i_0_9_lpi_1_dfm;
      COMP_i_0_10_lpi_1_dfm_5 <= COMP_i_0_10_lpi_1_dfm;
      COMP_i_0_11_lpi_1_dfm_5 <= COMP_i_0_11_lpi_1_dfm;
      COMP_i_0_12_lpi_1_dfm_5 <= COMP_i_0_12_lpi_1_dfm;
      COMP_i_0_13_lpi_1_dfm_5 <= COMP_i_0_13_lpi_1_dfm;
      COMP_i_0_14_lpi_1_dfm_5 <= COMP_i_0_14_lpi_1_dfm;
      COMP_i_0_15_lpi_1_dfm_5 <= COMP_i_0_15_lpi_1_dfm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_itm <= 1'b0;
    end
    else if ( and_235_itm & (~ exitL_exit_for_sva) & (~(exit_for_lpi_1_dfm_4 | lfst_exit_for_for_for_1_lpi_1_0_1))
        & core_wen ) begin
      reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_itm <= for_for_for_1_k_mux_itm[3];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_1_itm <=
          3'b0;
    end
    else if ( ((~(lfst_exit_for_for_for_1_lpi_1_1_1 & lfst_exit_for_for_1_lpi_2))
        | exitL_exit_for_sva | exit_for_lpi_1_dfm_4 | (~ lfst_exit_for_for_for_1_lpi_1_0_1))
        & core_wen ) begin
      reg_out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_4_1_1_itm <=
          for_for_for_1_k_mux_itm[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1 <= 1'b0;
    end
    else if ( core_wen & or_dcpl_18 ) begin
      out_stencil_operator_lo_out_stencil_operator_lo_conc_itm_1_0_1 <= MUX1HOT_s_1_3_2(for_for_for_1_for_q_0_lpi_2,
          (WX_if_1_acc_1_ncse[0]), pref_pref_pref_6_3_0_1_lpi_1_0_1, {and_dcpl_65
          , (or_75_nl) , (and_228_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_and_13_mdf_sva_6 <= 1'b0;
    end
    else if ( core_wen & (~((~((~((lfst_exit_for_for_for_1_lpi_1_dfm_1_st_4!=2'b00)
        | unequal_tmp_5)) & for_for_for_1_nor_dfs_5 & (~ lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1)
        & (for_for_row_6_0_lpi_1_dfm_9[6]))) & or_dcpl_13)) & main_stage_0_2 ) begin
      COMP_and_13_mdf_sva_6 <= COMP_and_13_mdf_sva_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      weight_buf_value_1_2_15_0_lpi_1 <= 16'b0;
      weight_buf_value_1_2_47_32_lpi_1 <= 16'b0;
    end
    else if ( weight_buf_value_and_cse ) begin
      weight_buf_value_1_2_15_0_lpi_1 <= weight_rsci_d_mxwt[15:0];
      weight_buf_value_1_2_47_32_lpi_1 <= weight_rsci_d_mxwt[31:16];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      weight_buf_value_0_1_15_0_lpi_1 <= 16'b0;
      weight_buf_value_0_1_47_32_lpi_1 <= 16'b0;
    end
    else if ( weight_buf_value_and_2_cse ) begin
      weight_buf_value_0_1_15_0_lpi_1 <= weight_rsci_d_mxwt[15:0];
      weight_buf_value_0_1_47_32_lpi_1 <= weight_rsci_d_mxwt[31:16];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      weight_buf_value_2_0_15_0_lpi_1 <= 16'b0;
      weight_buf_value_2_0_47_32_lpi_1 <= 16'b0;
    end
    else if ( weight_buf_value_and_4_cse ) begin
      weight_buf_value_2_0_15_0_lpi_1 <= weight_rsci_d_mxwt[15:0];
      weight_buf_value_2_0_47_32_lpi_1 <= weight_rsci_d_mxwt[31:16];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      weight_buf_value_0_2_15_0_lpi_1 <= 16'b0;
      weight_buf_value_0_2_47_32_lpi_1 <= 16'b0;
    end
    else if ( weight_buf_value_and_6_cse ) begin
      weight_buf_value_0_2_15_0_lpi_1 <= weight_rsci_d_mxwt[15:0];
      weight_buf_value_0_2_47_32_lpi_1 <= weight_rsci_d_mxwt[31:16];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      weight_buf_value_2_1_15_0_lpi_1 <= 16'b0;
      weight_buf_value_2_1_47_32_lpi_1 <= 16'b0;
    end
    else if ( weight_buf_value_and_8_cse ) begin
      weight_buf_value_2_1_15_0_lpi_1 <= weight_rsci_d_mxwt[15:0];
      weight_buf_value_2_1_47_32_lpi_1 <= weight_rsci_d_mxwt[31:16];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      weight_buf_value_1_0_15_0_lpi_1 <= 16'b0;
      weight_buf_value_1_0_47_32_lpi_1 <= 16'b0;
    end
    else if ( weight_buf_value_and_10_cse ) begin
      weight_buf_value_1_0_15_0_lpi_1 <= weight_rsci_d_mxwt[15:0];
      weight_buf_value_1_0_47_32_lpi_1 <= weight_rsci_d_mxwt[31:16];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      weight_buf_value_2_2_15_0_lpi_1 <= 16'b0;
      weight_buf_value_2_2_47_32_lpi_1 <= 16'b0;
    end
    else if ( weight_buf_value_and_12_cse ) begin
      weight_buf_value_2_2_15_0_lpi_1 <= weight_rsci_d_mxwt[15:0];
      weight_buf_value_2_2_47_32_lpi_1 <= weight_rsci_d_mxwt[31:16];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      weight_buf_value_0_0_15_0_lpi_1 <= 16'b0;
      weight_buf_value_0_0_47_32_lpi_1 <= 16'b0;
    end
    else if ( weight_buf_value_and_14_cse ) begin
      weight_buf_value_0_0_15_0_lpi_1 <= weight_rsci_d_mxwt[15:0];
      weight_buf_value_0_0_47_32_lpi_1 <= weight_rsci_d_mxwt[31:16];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      weight_buf_value_1_1_15_0_lpi_1 <= 16'b0;
      weight_buf_value_1_1_47_32_lpi_1 <= 16'b0;
    end
    else if ( weight_buf_value_and_16_cse ) begin
      weight_buf_value_1_1_15_0_lpi_1 <= weight_rsci_d_mxwt[15:0];
      weight_buf_value_1_1_47_32_lpi_1 <= weight_rsci_d_mxwt[31:16];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      WX_and_17_psp_1 <= 1'b0;
      WX_and_15_psp_1 <= 1'b0;
      WX_and_13_psp_1 <= 1'b0;
      WX_and_11_psp_1 <= 1'b0;
      WX_and_9_psp_1 <= 1'b0;
      WX_and_7_psp_1 <= 1'b0;
      WX_and_5_psp_1 <= 1'b0;
      WX_and_3_psp_1 <= 1'b0;
      WX_and_1_psp_1 <= 1'b0;
    end
    else if ( WX_and_19_cse ) begin
      WX_and_17_psp_1 <= WX_and_16_psp_mx0w0;
      WX_and_15_psp_1 <= WX_and_14_psp_mx0w0;
      WX_and_13_psp_1 <= WX_and_12_psp_mx0w0;
      WX_and_11_psp_1 <= WX_and_10_psp_mx0w0;
      WX_and_9_psp_1 <= WX_and_8_psp_mx0w0;
      WX_and_7_psp_1 <= WX_and_6_psp_mx0w0;
      WX_and_5_psp_1 <= WX_and_4_psp_mx0w0;
      WX_and_3_psp_1 <= WX_and_2_psp_mx0w0;
      WX_and_1_psp_1 <= WX_and_psp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      WX_if_1_and_stg_1_1_sva <= 1'b0;
      WX_if_1_and_stg_1_2_sva <= 1'b0;
      WX_if_1_and_stg_1_3_sva <= 1'b0;
      WX_if_1_and_stg_2_0_sva <= 1'b0;
      WX_if_1_and_stg_1_0_sva <= 1'b0;
    end
    else if ( WX_if_1_and_cse ) begin
      WX_if_1_and_stg_1_1_sva <= WX_if_1_and_stg_1_1_sva_mx0w0;
      WX_if_1_and_stg_1_2_sva <= WX_if_1_and_stg_1_2_sva_mx0w0;
      WX_if_1_and_stg_1_3_sva <= WX_if_1_and_stg_1_3_sva_mx0w0;
      WX_if_1_and_stg_2_0_sva <= WX_if_1_and_stg_2_0_sva_mx0w0;
      WX_if_1_and_stg_1_0_sva <= WX_if_1_and_stg_1_0_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_row_6_0_lpi_1_dfm_9 <= 7'b0;
    end
    else if ( core_wen & ((~((~((~ lfst_exit_for_for_for_1_lpi_1_0_1) | exitL_exit_COL_1_COMP_lpi_1
        | (~ lfst_exit_WX_1_lpi_1) | (~((WY_mux_6_tmp!=2'b00))))) | lfst_exit_for_for_for_1_lpi_1_1_1))
        | or_dcpl_13) ) begin
      for_for_row_6_0_lpi_1_dfm_9 <= for_for_row_6_0_lpi_1_dfm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      in_tmp_14_lpi_2 <= 16'b0;
    end
    else if ( core_wen & (((~ WX_unequal_tmp_5) & exitL_exit_COL_1_COMP_lpi_1_dfm_4
        & (~ for_for_for_1_or_cse) & main_stage_0_2) | and_119_rgt) & and_dcpl_38
        ) begin
      in_tmp_14_lpi_2 <= MUX_v_16_2_2((input_rsci_d_mxwt[239:224]), in_tmp_15_lpi_2,
          and_119_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      in_tmp_13_lpi_2 <= 16'b0;
      in_tmp_12_lpi_2 <= 16'b0;
      in_tmp_11_lpi_2 <= 16'b0;
      in_tmp_10_lpi_2 <= 16'b0;
      in_tmp_9_lpi_2 <= 16'b0;
      in_tmp_8_lpi_2 <= 16'b0;
      in_tmp_7_lpi_2 <= 16'b0;
      in_tmp_6_lpi_2 <= 16'b0;
      in_tmp_5_lpi_2 <= 16'b0;
      in_tmp_4_lpi_2 <= 16'b0;
      in_tmp_3_lpi_2 <= 16'b0;
      in_tmp_2_lpi_2 <= 16'b0;
      in_tmp_1_lpi_2 <= 16'b0;
    end
    else if ( in_tmp_and_1_cse ) begin
      in_tmp_13_lpi_2 <= in_tmp_14_lpi_1_dfm_1_mx0;
      in_tmp_12_lpi_2 <= in_tmp_13_lpi_1_dfm_1_mx0;
      in_tmp_11_lpi_2 <= in_tmp_12_lpi_1_dfm_1_mx0;
      in_tmp_10_lpi_2 <= in_tmp_11_lpi_1_dfm_1_mx0;
      in_tmp_9_lpi_2 <= in_tmp_10_lpi_1_dfm_1_mx0;
      in_tmp_8_lpi_2 <= in_tmp_9_lpi_1_dfm_1_mx0;
      in_tmp_7_lpi_2 <= in_tmp_8_lpi_1_dfm_1_mx0;
      in_tmp_6_lpi_2 <= in_tmp_7_lpi_1_dfm_1_mx0;
      in_tmp_5_lpi_2 <= in_tmp_6_lpi_1_dfm_1_mx0;
      in_tmp_4_lpi_2 <= in_tmp_5_lpi_1_dfm_1_mx0;
      in_tmp_3_lpi_2 <= in_tmp_4_lpi_1_dfm_1_mx0;
      in_tmp_2_lpi_2 <= in_tmp_3_lpi_1_dfm_1_mx0;
      in_tmp_1_lpi_2 <= in_tmp_2_lpi_1_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      in_tmp_15_lpi_2 <= 16'b0;
    end
    else if ( core_wen & ((asn_259 & (~(COMP_and_13_mdf_sva_5 | for_for_for_1_or_cse))
        & main_stage_0_2) | for_for_for_1_and_279_rgt) & or_tmp_19 & (~ exit_for_lpi_1_dfm_4)
        & (~ exitL_exit_for_sva) & lfst_exit_for_for_1_lpi_2 & and_dcpl_36 ) begin
      in_tmp_15_lpi_2 <= MUX_v_16_2_2((input_rsci_d_mxwt[239:224]), in_tmp_16_lpi_1_dfm_1,
          for_for_for_1_and_279_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pe_x_reg_13_lpi_2 <= 16'b0;
      pe_x_reg_12_lpi_2 <= 16'b0;
      pe_x_reg_11_lpi_2 <= 16'b0;
      pe_x_reg_10_lpi_2 <= 16'b0;
      pe_x_reg_9_lpi_2 <= 16'b0;
      pe_x_reg_8_lpi_2 <= 16'b0;
      pe_x_reg_7_lpi_2 <= 16'b0;
      pe_x_reg_6_lpi_2 <= 16'b0;
      pe_x_reg_5_lpi_2 <= 16'b0;
      pe_x_reg_4_lpi_2 <= 16'b0;
      pe_x_reg_3_lpi_2 <= 16'b0;
      pe_x_reg_2_lpi_2 <= 16'b0;
      pe_x_reg_1_lpi_2 <= 16'b0;
    end
    else if ( pe_x_reg_and_cse ) begin
      pe_x_reg_13_lpi_2 <= in_tmp_14_lpi_1_dfm_1_mx0;
      pe_x_reg_12_lpi_2 <= in_tmp_13_lpi_1_dfm_1_mx0;
      pe_x_reg_11_lpi_2 <= in_tmp_12_lpi_1_dfm_1_mx0;
      pe_x_reg_10_lpi_2 <= in_tmp_11_lpi_1_dfm_1_mx0;
      pe_x_reg_9_lpi_2 <= in_tmp_10_lpi_1_dfm_1_mx0;
      pe_x_reg_8_lpi_2 <= in_tmp_9_lpi_1_dfm_1_mx0;
      pe_x_reg_7_lpi_2 <= in_tmp_8_lpi_1_dfm_1_mx0;
      pe_x_reg_6_lpi_2 <= in_tmp_7_lpi_1_dfm_1_mx0;
      pe_x_reg_5_lpi_2 <= in_tmp_6_lpi_1_dfm_1_mx0;
      pe_x_reg_4_lpi_2 <= in_tmp_5_lpi_1_dfm_1_mx0;
      pe_x_reg_3_lpi_2 <= in_tmp_4_lpi_1_dfm_1_mx0;
      pe_x_reg_2_lpi_2 <= in_tmp_3_lpi_1_dfm_1_mx0;
      pe_x_reg_1_lpi_2 <= in_tmp_2_lpi_1_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_i_0_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & ((or_dcpl_9 & (~ lfst_exit_for_for_for_1_lpi_1_0_1) & (for_for_for_1_acc_1_tmp[4])
        & for_for_for_1_for_q_0_lpi_2 & for_for_for_1_nand_2_tmp) | or_71_cse) )
        begin
      COMP_i_0_1_lpi_1_dfm_5 <= MUX_s_1_2_2(COMP_i_0_1_lpi_1_dfm, (for_for_acc_1_tmp[6]),
          and_dcpl_65);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      in_tmp_16_lpi_2 <= 16'b0;
      pe_x_reg_0_lpi_2 <= 16'b0;
    end
    else if ( in_tmp_and_14_cse ) begin
      in_tmp_16_lpi_2 <= in_tmp_16_lpi_1_dfm_1;
      pe_x_reg_0_lpi_2 <= pe_x_reg_0_lpi_1_dfm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_for_1_nor_dfs_6 <= 1'b0;
      unequal_tmp_6 <= 1'b0;
      lfst_exit_for_for_for_1_lpi_1_dfm_9_1_1 <= 1'b0;
    end
    else if ( for_for_for_1_and_300_cse ) begin
      for_for_for_1_nor_dfs_6 <= for_for_for_1_nor_dfs_5;
      unequal_tmp_6 <= unequal_tmp_5;
      lfst_exit_for_for_for_1_lpi_1_dfm_9_1_1 <= slc_lfst_exit_for_for_for_1_1_1_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      for_for_row_6_0_lpi_1_dfm_6_6_1 <= 1'b0;
    end
    else if ( core_wen & (mux_159_nl) & main_stage_0_2 ) begin
      for_for_row_6_0_lpi_1_dfm_6_6_1 <= MUX_s_1_2_2((for_for_row_6_0_lpi_1_dfm_9[6]),
          COMP_i_0_1_lpi_1_dfm_5, lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_and_13_mdf_sva_5 <= 1'b0;
    end
    else if ( core_wen & (mux_160_nl) ) begin
      COMP_and_13_mdf_sva_5 <= COMP_and_13_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      WX_if_1_acc_decb_sva_3_1 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_61) ) begin
      WX_if_1_acc_decb_sva_3_1 <= WX_if_1_acc_decb_sva_3_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pref_pref_pref_6_3_0_1_lpi_1_3_1_1 <= 3'b0;
      pref_pref_pref_6_3_0_1_lpi_1_0_1 <= 1'b0;
    end
    else if ( COL_and_cse ) begin
      pref_pref_pref_6_3_0_1_lpi_1_3_1_1 <= WX_if_1_acc_decb_sva_3_1_mx0w0;
      pref_pref_pref_6_3_0_1_lpi_1_0_1 <= WX_if_1_acc_1_ncse[0];
    end
  end
  assign for_for_for_1_mux1h_196_nl = MUX1HOT_s_1_4_2((for_for_row_6_0_lpi_1_dfm[6]),
      (WY_mux_3_cse[1]), (~ exit_for_for_for_1_lpi_1_dfm_1), lfst_exit_for_for_for_1_lpi_1_dfm_1,
      {for_for_for_1_and_3_cse , for_for_for_1_and_4_m1c , for_for_for_1_and_96_cse
      , for_for_for_1_equal_tmp_1});
  assign for_for_for_1_mux1h_193_nl = MUX1HOT_s_1_3_2((for_for_row_6_0_lpi_1_dfm[6]),
      (WY_mux_3_cse[0]), lfst_exit_for_for_for_1_lpi_1_dfm_0, {for_for_for_1_and_3_cse
      , for_for_for_1_and_4_m1c , for_for_for_1_equal_tmp_1});
  assign or_68_nl = (~ exitL_exit_COL_1_COMP_lpi_1_dfm_4) | WX_unequal_tmp_5;
  assign and_233_nl = ((for_for_row_6_0_lpi_3[5:0]!=6'b000000)) & lfst_exit_for_lpi_1_dfm;
  assign WY_not_10_nl = ~ exit_WY_lpi_1_dfm_2;
  assign WY_WY_and_2_nl = MUX_v_4_2_2(4'b0000, for_for_for_1_k_4_0_lpi_1_3_0_1, (WY_not_10_nl));
  assign nor_60_nl = ~((~ COMP_and_13_tmp) | WX_acc_tmp_1 | WY_acc_tmp_1);
  assign nor_61_nl = ~(lfst_exit_for_for_for_1_lpi_1_0_1 | (~ for_for_for_1_for_q_0_lpi_2));
  assign or_170_nl = (~ lfst_exit_for_for_for_1_lpi_1_1_1) | (~ lfst_exit_for_for_1_lpi_2)
      | exit_for_lpi_1_dfm_4 | exitL_exit_for_sva;
  assign mux_201_nl = MUX_s_1_2_2((nor_61_nl), (nor_60_nl), or_170_nl);
  assign WY_WY_and_3_nl = for_for_for_1_for_q_0_lpi_2 & (~ exit_WY_lpi_1_dfm_2);
  assign and_55_nl = (~ for_for_for_1_for_q_0_lpi_2) & (for_for_for_1_acc_1_tmp[4]);
  assign and_241_nl = (((for_for_row_6_0_lpi_1_dfm[6]) & for_for_for_1_and_3_cse)
      | for_for_for_1_and_4_m1c) & exit_WX_lpi_1_dfm_1;
  assign mux_203_nl = MUX_v_2_2_2(WY_wy_1_0_lpi_1_dfm, WY_wy_1_0_sva_1, and_241_nl);
  assign nor_64_nl = ~(((~ (for_for_acc_1_tmp[6])) & for_for_for_1_and_95_cse) |
      ((~ (for_for_row_6_0_lpi_1_dfm[6])) & for_for_for_1_and_3_cse));
  assign for_for_for_1_nand_nl = ~(for_for_for_1_equal_tmp & (~((~ exit_for_for_for_1_lpi_1_dfm_1)
      & for_for_for_1_and_2_m1c)));
  assign for_for_for_1_and_nl = exit_for_for_lpi_1_dfm_5 & for_for_for_1_equal_tmp;
  assign for_for_for_1_and_166_nl = exit_for_for_for_1_lpi_1_dfm_1 & for_for_for_1_and_2_m1c;
  assign and_232_nl = and_dcpl_65 & (~ lfst_exit_for_for_for_1_lpi_1_0_1) & (for_for_for_1_acc_1_tmp[4])
      & for_for_for_1_for_q_0_lpi_2 & (for_for_acc_1_tmp[6]);
  assign and_59_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_0_31_0_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign mux_204_nl = MUX_s_1_2_2(not_tmp_131, or_tmp_84, main_stage_0_3);
  assign nand_10_nl = ~(lfst_exit_for_for_1_lpi_1_dfm_1 & (~ (mux_204_nl)));
  assign or_202_nl = (~ lfst_exit_for_for_1_lpi_2) | exitL_exit_for_sva | exit_for_lpi_1_dfm_4
      | not_tmp_131;
  assign mux_205_nl = MUX_s_1_2_2((or_202_nl), or_tmp_84, main_stage_0_3);
  assign mux_206_nl = MUX_s_1_2_2((mux_205_nl), (nand_10_nl), main_stage_0_2);
  assign and_259_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_7_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_316_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_207_nl = MUX_s_1_2_2(nor_317_cse, (nor_316_nl), COMP_and_13_mdf_sva_6);
  assign nor_315_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_207_nl));
  assign mux_208_nl = MUX_s_1_2_2((nor_315_nl), (and_259_nl), unequal_tmp_6);
  assign and_264_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_7_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_313_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_209_nl = MUX_s_1_2_2(nor_317_cse, (nor_313_nl), COMP_and_13_mdf_sva_6);
  assign nor_312_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_209_nl));
  assign mux_210_nl = MUX_s_1_2_2((nor_312_nl), (and_264_nl), unequal_tmp_6);
  assign and_269_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_6_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_310_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_15_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_211_nl = MUX_s_1_2_2(nor_317_cse, (nor_310_nl), COMP_and_13_mdf_sva_6);
  assign nor_309_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_211_nl));
  assign mux_212_nl = MUX_s_1_2_2((nor_309_nl), (and_269_nl), unequal_tmp_6);
  assign and_274_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_6_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_307_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_15_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_213_nl = MUX_s_1_2_2(nor_317_cse, (nor_307_nl), COMP_and_13_mdf_sva_6);
  assign nor_306_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_213_nl));
  assign mux_214_nl = MUX_s_1_2_2((nor_306_nl), (and_274_nl), unequal_tmp_6);
  assign and_279_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_5_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_304_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_14_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_215_nl = MUX_s_1_2_2(nor_317_cse, (nor_304_nl), COMP_and_13_mdf_sva_6);
  assign nor_303_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_215_nl));
  assign mux_216_nl = MUX_s_1_2_2((nor_303_nl), (and_279_nl), unequal_tmp_6);
  assign and_284_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_4_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_301_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_14_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_217_nl = MUX_s_1_2_2(nor_317_cse, (nor_301_nl), COMP_and_13_mdf_sva_6);
  assign nor_300_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_217_nl));
  assign mux_218_nl = MUX_s_1_2_2((nor_300_nl), (and_284_nl), unequal_tmp_6);
  assign and_289_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_4_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_298_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_13_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_219_nl = MUX_s_1_2_2(nor_317_cse, (nor_298_nl), COMP_and_13_mdf_sva_6);
  assign nor_297_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_219_nl));
  assign mux_220_nl = MUX_s_1_2_2((nor_297_nl), (and_289_nl), unequal_tmp_6);
  assign and_294_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_3_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_295_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_13_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_221_nl = MUX_s_1_2_2(nor_317_cse, (nor_295_nl), COMP_and_13_mdf_sva_6);
  assign nor_294_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_221_nl));
  assign mux_222_nl = MUX_s_1_2_2((nor_294_nl), (and_294_nl), unequal_tmp_6);
  assign and_299_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_3_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_292_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_12_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_223_nl = MUX_s_1_2_2(nor_317_cse, (nor_292_nl), COMP_and_13_mdf_sva_6);
  assign nor_291_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_223_nl));
  assign mux_224_nl = MUX_s_1_2_2((nor_291_nl), (and_299_nl), unequal_tmp_6);
  assign and_304_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_289_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_12_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_225_nl = MUX_s_1_2_2(nor_317_cse, (nor_289_nl), COMP_and_13_mdf_sva_6);
  assign nor_288_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_225_nl));
  assign mux_226_nl = MUX_s_1_2_2((nor_288_nl), (and_304_nl), unequal_tmp_6);
  assign and_309_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_286_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_11_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_227_nl = MUX_s_1_2_2(nor_317_cse, (nor_286_nl), COMP_and_13_mdf_sva_6);
  assign nor_285_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_227_nl));
  assign mux_228_nl = MUX_s_1_2_2((nor_285_nl), (and_309_nl), unequal_tmp_6);
  assign and_314_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_15_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_283_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_11_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_229_nl = MUX_s_1_2_2(nor_317_cse, (nor_283_nl), COMP_and_13_mdf_sva_6);
  assign nor_282_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_229_nl));
  assign mux_230_nl = MUX_s_1_2_2((nor_282_nl), (and_314_nl), unequal_tmp_6);
  assign and_319_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_15_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_280_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_10_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_231_nl = MUX_s_1_2_2(nor_317_cse, (nor_280_nl), COMP_and_13_mdf_sva_6);
  assign nor_279_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_231_nl));
  assign mux_232_nl = MUX_s_1_2_2((nor_279_nl), (and_319_nl), unequal_tmp_6);
  assign and_324_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_14_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_277_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_10_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_233_nl = MUX_s_1_2_2(nor_317_cse, (nor_277_nl), COMP_and_13_mdf_sva_6);
  assign nor_276_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_233_nl));
  assign mux_234_nl = MUX_s_1_2_2((nor_276_nl), (and_324_nl), unequal_tmp_6);
  assign and_329_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_13_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_274_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_9_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_235_nl = MUX_s_1_2_2(nor_317_cse, (nor_274_nl), COMP_and_13_mdf_sva_6);
  assign nor_273_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_235_nl));
  assign mux_236_nl = MUX_s_1_2_2((nor_273_nl), (and_329_nl), unequal_tmp_6);
  assign and_334_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_13_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_271_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_9_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_237_nl = MUX_s_1_2_2(nor_317_cse, (nor_271_nl), COMP_and_13_mdf_sva_6);
  assign nor_270_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_237_nl));
  assign mux_238_nl = MUX_s_1_2_2((nor_270_nl), (and_334_nl), unequal_tmp_6);
  assign and_339_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_12_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_268_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_8_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_239_nl = MUX_s_1_2_2(nor_317_cse, (nor_268_nl), COMP_and_13_mdf_sva_6);
  assign nor_267_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_239_nl));
  assign mux_240_nl = MUX_s_1_2_2((nor_267_nl), (and_339_nl), unequal_tmp_6);
  assign and_344_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_12_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_265_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_8_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_241_nl = MUX_s_1_2_2(nor_317_cse, (nor_265_nl), COMP_and_13_mdf_sva_6);
  assign nor_264_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_241_nl));
  assign mux_242_nl = MUX_s_1_2_2((nor_264_nl), (and_344_nl), unequal_tmp_6);
  assign and_349_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_11_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_262_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_7_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_243_nl = MUX_s_1_2_2(nor_317_cse, (nor_262_nl), COMP_and_13_mdf_sva_6);
  assign nor_261_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_243_nl));
  assign mux_244_nl = MUX_s_1_2_2((nor_261_nl), (and_349_nl), unequal_tmp_6);
  assign and_354_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_11_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_259_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_7_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_245_nl = MUX_s_1_2_2(nor_317_cse, (nor_259_nl), COMP_and_13_mdf_sva_6);
  assign nor_258_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_245_nl));
  assign mux_246_nl = MUX_s_1_2_2((nor_258_nl), (and_354_nl), unequal_tmp_6);
  assign and_359_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_2_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_256_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_6_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_247_nl = MUX_s_1_2_2(nor_317_cse, (nor_256_nl), COMP_and_13_mdf_sva_6);
  assign nor_255_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_247_nl));
  assign mux_248_nl = MUX_s_1_2_2((nor_255_nl), (and_359_nl), unequal_tmp_6);
  assign and_364_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_2_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_253_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_6_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_249_nl = MUX_s_1_2_2(nor_317_cse, (nor_253_nl), COMP_and_13_mdf_sva_6);
  assign nor_252_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_249_nl));
  assign mux_250_nl = MUX_s_1_2_2((nor_252_nl), (and_364_nl), unequal_tmp_6);
  assign and_369_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_1_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_250_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_5_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_251_nl = MUX_s_1_2_2(nor_317_cse, (nor_250_nl), COMP_and_13_mdf_sva_6);
  assign nor_249_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_251_nl));
  assign mux_252_nl = MUX_s_1_2_2((nor_249_nl), (and_369_nl), unequal_tmp_6);
  assign and_374_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_1_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_247_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_5_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_253_nl = MUX_s_1_2_2(nor_317_cse, (nor_247_nl), COMP_and_13_mdf_sva_6);
  assign nor_246_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_253_nl));
  assign mux_254_nl = MUX_s_1_2_2((nor_246_nl), (and_374_nl), unequal_tmp_6);
  assign and_379_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_10_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_244_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_4_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_255_nl = MUX_s_1_2_2(nor_317_cse, (nor_244_nl), COMP_and_13_mdf_sva_6);
  assign nor_243_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_255_nl));
  assign mux_256_nl = MUX_s_1_2_2((nor_243_nl), (and_379_nl), unequal_tmp_6);
  assign and_384_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_10_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_241_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_4_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_257_nl = MUX_s_1_2_2(nor_317_cse, (nor_241_nl), COMP_and_13_mdf_sva_6);
  assign nor_240_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_257_nl));
  assign mux_258_nl = MUX_s_1_2_2((nor_240_nl), (and_384_nl), unequal_tmp_6);
  assign and_389_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_9_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_238_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_3_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_259_nl = MUX_s_1_2_2(nor_317_cse, (nor_238_nl), COMP_and_13_mdf_sva_6);
  assign nor_237_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_259_nl));
  assign mux_260_nl = MUX_s_1_2_2((nor_237_nl), (and_389_nl), unequal_tmp_6);
  assign and_394_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_9_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_235_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_3_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_261_nl = MUX_s_1_2_2(nor_317_cse, (nor_235_nl), COMP_and_13_mdf_sva_6);
  assign nor_234_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_261_nl));
  assign mux_262_nl = MUX_s_1_2_2((nor_234_nl), (and_394_nl), unequal_tmp_6);
  assign and_399_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_8_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_232_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_2_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_263_nl = MUX_s_1_2_2(nor_317_cse, (nor_232_nl), COMP_and_13_mdf_sva_6);
  assign nor_231_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_263_nl));
  assign mux_264_nl = MUX_s_1_2_2((nor_231_nl), (and_399_nl), unequal_tmp_6);
  assign and_404_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_8_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_229_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_2_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_265_nl = MUX_s_1_2_2(nor_317_cse, (nor_229_nl), COMP_and_13_mdf_sva_6);
  assign nor_228_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_265_nl));
  assign mux_266_nl = MUX_s_1_2_2((nor_228_nl), (and_404_nl), unequal_tmp_6);
  assign and_409_nl = COMP_and_13_mdf_sva_6 & (COMP_i_0_5_lpi_1_dfm_6 | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_226_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | (~ COMP_i_0_1_lpi_1_dfm_6)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_267_nl = MUX_s_1_2_2(nor_317_cse, (nor_226_nl), COMP_and_13_mdf_sva_6);
  assign nor_225_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_267_nl));
  assign mux_268_nl = MUX_s_1_2_2((nor_225_nl), (and_409_nl), unequal_tmp_6);
  assign and_414_nl = COMP_and_13_mdf_sva_6 & ((~ COMP_i_0_14_lpi_1_dfm_6) | (~ exit_for_for_for_1_lpi_1_dfm_1_st_4)
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign nor_223_nl = ~((~ exit_for_for_for_1_lpi_1_dfm_1_st_4) | COMP_i_0_1_lpi_1_dfm_6
      | (~ lfst_exit_for_for_1_lpi_1_dfm_4) | (~ main_stage_0_4) | for_for_for_1_nor_dfs_7
      | for_for_for_1_equal_tmp_11 | for_for_for_1_equal_tmp_13);
  assign mux_269_nl = MUX_s_1_2_2(nor_317_cse, (nor_223_nl), COMP_and_13_mdf_sva_6);
  assign nor_222_nl = ~((~ for_for_row_6_0_lpi_1_dfm_6_6_1) | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_5!=2'b00)
      | lfst_exit_for_for_for_1_lpi_1_dfm_st_2_1_1 | (mux_269_nl));
  assign mux_270_nl = MUX_s_1_2_2((nor_222_nl), (and_414_nl), unequal_tmp_6);
  assign and_89_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_15_31_0_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_88_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_15_63_32_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_87_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_14_31_0_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_86_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_14_63_32_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_85_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_13_31_0_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_84_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_13_63_32_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_83_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_12_31_0_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_82_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_12_63_32_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_81_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_11_31_0_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_80_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_11_63_32_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_79_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_10_31_0_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_78_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_10_63_32_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_61_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_1_31_0_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_60_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_1_63_32_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign and_58_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000, out_tmp_value_0_63_32_lpi_1_dfm_mx0w0,
      for_for_row_6_0_lpi_1_dfm_6_6_1);
  assign nor_321_nl = ~(COMP_i_0_1_lpi_1_dfm_5 | and_741_tmp);
  assign and_751_nl = COMP_i_0_1_lpi_1_dfm_5 & (~ and_741_tmp);
  assign mux1h_nl = MUX1HOT_v_16_3_2(weight_buf_value_2_2_15_0_lpi_1, weight_buf_value_2_2_47_32_lpi_1,
      mux_414_cse, {(nor_321_nl) , (and_751_nl) , and_741_tmp});
  assign nor_322_nl = ~(COMP_i_0_1_lpi_1_dfm_5 | and_742_tmp);
  assign and_753_nl = COMP_i_0_1_lpi_1_dfm_5 & (~ and_742_tmp);
  assign mux1h_38_nl = MUX1HOT_v_16_3_2(weight_buf_value_2_1_15_0_lpi_1, weight_buf_value_2_1_47_32_lpi_1,
      mux_414_cse, {(nor_322_nl) , (and_753_nl) , and_742_tmp});
  assign nor_323_nl = ~(COMP_i_0_1_lpi_1_dfm_5 | and_743_tmp);
  assign and_755_nl = COMP_i_0_1_lpi_1_dfm_5 & (~ and_743_tmp);
  assign mux1h_39_nl = MUX1HOT_v_16_3_2(weight_buf_value_2_0_15_0_lpi_1, weight_buf_value_2_0_47_32_lpi_1,
      mux_414_cse, {(nor_323_nl) , (and_755_nl) , and_743_tmp});
  assign nor_324_nl = ~(COMP_i_0_1_lpi_1_dfm_5 | and_744_tmp);
  assign and_757_nl = COMP_i_0_1_lpi_1_dfm_5 & (~ and_744_tmp);
  assign mux1h_40_nl = MUX1HOT_v_16_3_2(weight_buf_value_1_2_15_0_lpi_1, weight_buf_value_1_2_47_32_lpi_1,
      mux_414_cse, {(nor_324_nl) , (and_757_nl) , and_744_tmp});
  assign nor_325_nl = ~(COMP_i_0_1_lpi_1_dfm_5 | and_745_tmp);
  assign and_759_nl = COMP_i_0_1_lpi_1_dfm_5 & (~ and_745_tmp);
  assign mux1h_41_nl = MUX1HOT_v_16_3_2(weight_buf_value_1_1_15_0_lpi_1, weight_buf_value_1_1_47_32_lpi_1,
      mux_414_cse, {(nor_325_nl) , (and_759_nl) , and_745_tmp});
  assign nor_326_nl = ~(COMP_i_0_1_lpi_1_dfm_5 | and_746_tmp);
  assign and_761_nl = COMP_i_0_1_lpi_1_dfm_5 & (~ and_746_tmp);
  assign mux1h_42_nl = MUX1HOT_v_16_3_2(weight_buf_value_1_0_15_0_lpi_1, weight_buf_value_1_0_47_32_lpi_1,
      mux_414_cse, {(nor_326_nl) , (and_761_nl) , and_746_tmp});
  assign nor_327_nl = ~(COMP_i_0_1_lpi_1_dfm_5 | and_747_tmp);
  assign and_763_nl = COMP_i_0_1_lpi_1_dfm_5 & (~ and_747_tmp);
  assign mux1h_43_nl = MUX1HOT_v_16_3_2(weight_buf_value_0_2_15_0_lpi_1, weight_buf_value_0_2_47_32_lpi_1,
      mux_414_cse, {(nor_327_nl) , (and_763_nl) , and_747_tmp});
  assign nor_328_nl = ~(COMP_i_0_1_lpi_1_dfm_5 | and_748_tmp);
  assign and_765_nl = COMP_i_0_1_lpi_1_dfm_5 & (~ and_748_tmp);
  assign mux1h_44_nl = MUX1HOT_v_16_3_2(weight_buf_value_0_1_15_0_lpi_1, weight_buf_value_0_1_47_32_lpi_1,
      mux_414_cse, {(nor_328_nl) , (and_765_nl) , and_748_tmp});
  assign nor_329_nl = ~(COMP_i_0_1_lpi_1_dfm_5 | and_749_tmp);
  assign and_767_nl = COMP_i_0_1_lpi_1_dfm_5 & (~ and_749_tmp);
  assign mux1h_45_nl = MUX1HOT_v_16_3_2(weight_buf_value_0_0_15_0_lpi_1, weight_buf_value_0_0_47_32_lpi_1,
      mux_414_cse, {(nor_329_nl) , (and_767_nl) , and_749_tmp});
  assign or_75_nl = nor_41_cse | or_dcpl_7 | (~ lfst_exit_for_for_1_lpi_2);
  assign and_228_nl = lfst_exit_for_lpi_1_dfm & lfst_exit_for_for_1_lpi_2 & (~ lfst_exit_for_for_for_1_lpi_1_1_1)
      & and_dcpl_59;
  assign nor_45_nl = ~(slc_lfst_exit_for_for_for_1_1_1_itm_4 | lfst_exit_for_for_for_1_lpi_1_dfm_st_1_0
      | (~ for_for_for_1_equal_tmp_2) | (~ lfst_exit_for_for_1_lpi_2) | exitL_exit_for_sva
      | exit_for_lpi_1_dfm_4);
  assign nor_46_nl = ~((~ for_for_for_1_nor_dfs_5) | unequal_tmp_5 | (lfst_exit_for_for_for_1_lpi_1_dfm_1_st_4!=2'b00));
  assign mux_159_nl = MUX_s_1_2_2((nor_46_nl), (nor_45_nl), lfst_exit_for_for_for_1_lpi_1_dfm_st_1_1);
  assign nor_44_nl = ~((WY_mux_6_tmp[0]) | (~ (for_for_row_6_0_lpi_3[6])) | (WY_mux_6_tmp[1])
      | and_235_itm | exitL_exit_for_sva | exit_for_lpi_1_dfm_4);
  assign mux_160_nl = MUX_s_1_2_2((nor_44_nl), or_dcpl_15, for_for_for_1_nand_2_tmp);

  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function [31:0] MUX1HOT_v_32_4_2;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [3:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    MUX1HOT_v_32_4_2 = result;
  end
  endfunction


  function [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function [15:0] MUX_v_16_9_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [3:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      default : begin
        result = input_8;
      end
    endcase
    MUX_v_16_9_2 = result;
  end
  endfunction


  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [31:0] MUX_v_32_16_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [3:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_32_16_2 = result;
  end
  endfunction


  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function [6:0] signext_7_1;
    input [0:0] vector;
  begin
    signext_7_1= {{6{vector[0]}}, vector};
  end
  endfunction


  function [1023:0] writeslice_1024_5_32;
    input [1023:0] vector;
    input [31:0] slice;
    input [4:0] index;
    input esize;
    integer esize;
    input offs;
    integer offs;
    integer i;
    reg [1023:0] rvalue;
  begin
    rvalue = vector;
    for (i = 0; i < 32; i = i+1)
      rvalue[index * esize + offs + i] = slice[i];
    writeslice_1024_5_32 = rvalue;
  end
  endfunction


  function  [16:0] conv_u2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2s_16_17 =  {1'b0, vector};
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function  [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function  [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, dout_0_rsc_req_vz, dout_0_rsc_rls_lz,
      dout_1_rsc_req_vz, dout_1_rsc_rls_lz, dout_2_rsc_req_vz, dout_2_rsc_rls_lz,
      dout_3_rsc_req_vz, dout_3_rsc_rls_lz, dout_4_rsc_req_vz, dout_4_rsc_rls_lz,
      dout_5_rsc_req_vz, dout_5_rsc_rls_lz, dout_6_rsc_req_vz, dout_6_rsc_rls_lz,
      dout_7_rsc_req_vz, dout_7_rsc_rls_lz, dout_8_rsc_req_vz, dout_8_rsc_rls_lz,
      dout_9_rsc_req_vz, dout_9_rsc_rls_lz, dout_10_rsc_req_vz, dout_10_rsc_rls_lz,
      dout_11_rsc_req_vz, dout_11_rsc_rls_lz, dout_12_rsc_req_vz, dout_12_rsc_rls_lz,
      dout_13_rsc_req_vz, dout_13_rsc_rls_lz, dout_14_rsc_req_vz, dout_14_rsc_rls_lz,
      dout_15_rsc_req_vz, dout_15_rsc_rls_lz, dout_0_rsci_addra_d, dout_0_rsci_addrb_d,
      dout_0_rsci_dinb_d, dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d, dout_1_rsci_addra_d,
      dout_1_rsci_addrb_d, dout_1_rsci_dinb_d, dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_2_rsci_addra_d, dout_2_rsci_addrb_d, dout_2_rsci_dinb_d, dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_3_rsci_addra_d, dout_3_rsci_addrb_d, dout_3_rsci_dinb_d, dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_4_rsci_addra_d, dout_4_rsci_addrb_d, dout_4_rsci_dinb_d, dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_5_rsci_addra_d, dout_5_rsci_addrb_d, dout_5_rsci_dinb_d, dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_6_rsci_addra_d, dout_6_rsci_addrb_d, dout_6_rsci_dinb_d, dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_7_rsci_addra_d, dout_7_rsci_addrb_d, dout_7_rsci_dinb_d, dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_8_rsci_addra_d, dout_8_rsci_addrb_d, dout_8_rsci_dinb_d, dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_9_rsci_addra_d, dout_9_rsci_addrb_d, dout_9_rsci_dinb_d, dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_10_rsci_addra_d, dout_10_rsci_addrb_d, dout_10_rsci_dinb_d, dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_11_rsci_addra_d, dout_11_rsci_addrb_d, dout_11_rsci_dinb_d, dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_12_rsci_addra_d, dout_12_rsci_addrb_d, dout_12_rsci_dinb_d, dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_13_rsci_addra_d, dout_13_rsci_addrb_d, dout_13_rsci_dinb_d, dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_14_rsci_addra_d, dout_14_rsci_addrb_d, dout_14_rsci_dinb_d, dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d,
      dout_15_rsci_addra_d, dout_15_rsci_addrb_d, dout_15_rsci_dinb_d, dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d
);
  input clk;
  input rst;
  input [1023:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  input dout_0_rsc_req_vz;
  output dout_0_rsc_rls_lz;
  input dout_1_rsc_req_vz;
  output dout_1_rsc_rls_lz;
  input dout_2_rsc_req_vz;
  output dout_2_rsc_rls_lz;
  input dout_3_rsc_req_vz;
  output dout_3_rsc_rls_lz;
  input dout_4_rsc_req_vz;
  output dout_4_rsc_rls_lz;
  input dout_5_rsc_req_vz;
  output dout_5_rsc_rls_lz;
  input dout_6_rsc_req_vz;
  output dout_6_rsc_rls_lz;
  input dout_7_rsc_req_vz;
  output dout_7_rsc_rls_lz;
  input dout_8_rsc_req_vz;
  output dout_8_rsc_rls_lz;
  input dout_9_rsc_req_vz;
  output dout_9_rsc_rls_lz;
  input dout_10_rsc_req_vz;
  output dout_10_rsc_rls_lz;
  input dout_11_rsc_req_vz;
  output dout_11_rsc_rls_lz;
  input dout_12_rsc_req_vz;
  output dout_12_rsc_rls_lz;
  input dout_13_rsc_req_vz;
  output dout_13_rsc_rls_lz;
  input dout_14_rsc_req_vz;
  output dout_14_rsc_rls_lz;
  input dout_15_rsc_req_vz;
  output dout_15_rsc_rls_lz;
  output [7:0] dout_0_rsci_addra_d;
  output [7:0] dout_0_rsci_addrb_d;
  output [63:0] dout_0_rsci_dinb_d;
  output dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_1_rsci_addra_d;
  output [7:0] dout_1_rsci_addrb_d;
  output [63:0] dout_1_rsci_dinb_d;
  output dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_2_rsci_addra_d;
  output [7:0] dout_2_rsci_addrb_d;
  output [63:0] dout_2_rsci_dinb_d;
  output dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_3_rsci_addra_d;
  output [7:0] dout_3_rsci_addrb_d;
  output [63:0] dout_3_rsci_dinb_d;
  output dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_4_rsci_addra_d;
  output [7:0] dout_4_rsci_addrb_d;
  output [63:0] dout_4_rsci_dinb_d;
  output dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_5_rsci_addra_d;
  output [7:0] dout_5_rsci_addrb_d;
  output [63:0] dout_5_rsci_dinb_d;
  output dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_6_rsci_addra_d;
  output [7:0] dout_6_rsci_addrb_d;
  output [63:0] dout_6_rsci_dinb_d;
  output dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_7_rsci_addra_d;
  output [7:0] dout_7_rsci_addrb_d;
  output [63:0] dout_7_rsci_dinb_d;
  output dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_8_rsci_addra_d;
  output [7:0] dout_8_rsci_addrb_d;
  output [63:0] dout_8_rsci_dinb_d;
  output dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_9_rsci_addra_d;
  output [7:0] dout_9_rsci_addrb_d;
  output [63:0] dout_9_rsci_dinb_d;
  output dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_10_rsci_addra_d;
  output [7:0] dout_10_rsci_addrb_d;
  output [63:0] dout_10_rsci_dinb_d;
  output dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_11_rsci_addra_d;
  output [7:0] dout_11_rsci_addrb_d;
  output [63:0] dout_11_rsci_dinb_d;
  output dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_12_rsci_addra_d;
  output [7:0] dout_12_rsci_addrb_d;
  output [63:0] dout_12_rsci_dinb_d;
  output dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_13_rsci_addra_d;
  output [7:0] dout_13_rsci_addrb_d;
  output [63:0] dout_13_rsci_dinb_d;
  output dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_14_rsci_addra_d;
  output [7:0] dout_14_rsci_addrb_d;
  output [63:0] dout_14_rsci_dinb_d;
  output dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  output [7:0] dout_15_rsci_addra_d;
  output [7:0] dout_15_rsci_addrb_d;
  output [63:0] dout_15_rsci_dinb_d;
  output dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;


  // Interconnect Declarations
  wire core_wen;
  wire din_rsci_wen_comp;
  wire [1023:0] din_rsci_d_mxwt;
  wire core_wten;
  wire dout_15_rsc_req_obj_wen_comp;
  wire dout_14_rsc_req_obj_wen_comp;
  wire dout_13_rsc_req_obj_wen_comp;
  wire dout_12_rsc_req_obj_wen_comp;
  wire dout_11_rsc_req_obj_wen_comp;
  wire dout_10_rsc_req_obj_wen_comp;
  wire dout_9_rsc_req_obj_wen_comp;
  wire dout_8_rsc_req_obj_wen_comp;
  wire dout_7_rsc_req_obj_wen_comp;
  wire dout_6_rsc_req_obj_wen_comp;
  wire dout_5_rsc_req_obj_wen_comp;
  wire dout_4_rsc_req_obj_wen_comp;
  wire dout_3_rsc_req_obj_wen_comp;
  wire dout_2_rsc_req_obj_wen_comp;
  wire dout_1_rsc_req_obj_wen_comp;
  wire dout_0_rsc_req_obj_wen_comp;
  wire [1:0] fsm_output;
  wire [6:0] WRITE_acc_17_tmp;
  wire [7:0] nl_WRITE_acc_17_tmp;
  reg exitL_exit_for_sva;
  reg exit_for_lpi_1_dfm_2;
  reg [1:0] for_k_idx_2_0_lpi_1_dfm_1_1_0_1;
  reg [5:0] WRITE_y_idx_6_0_lpi_1_dfm_2_5_0_2;
  wire [2:0] for_k_idx_2_0_sva_1;
  wire [3:0] nl_for_k_idx_2_0_sva_1;
  reg reg_dout_15_rsc_req_obj_oswt_cse;
  reg reg_dout_0_rsc_rls_obj_ld_core_psct_cse;
  reg reg_din_rsci_ld_core_psct_cse;
  wire for_and_cse;
  wire nand_1_cse;
  wire dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire [1:0] for_k_idx_2_0_lpi_1_dfm_1_0;
  wire [5:0] WRITE_y_idx_6_0_lpi_1_dfm_5_0;
  wire exit_for_lpi_1_dfm_2_mx0w0;
  wire WRITE_y_idx_and_cse;

  wire[0:0] nor_nl;
  wire[0:0] for_not_7_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_inst_dout_0_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_inst_dout_0_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_inst_dout_1_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_inst_dout_1_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_inst_dout_2_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_inst_dout_2_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_inst_dout_3_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_inst_dout_3_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_inst_dout_4_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_inst_dout_4_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_inst_dout_5_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_inst_dout_5_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_inst_dout_6_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_inst_dout_6_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_inst_dout_7_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_inst_dout_7_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_inst_dout_8_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_inst_dout_8_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_inst_dout_9_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_inst_dout_9_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_inst_dout_10_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_inst_dout_10_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_inst_dout_11_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_inst_dout_11_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_inst_dout_12_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_inst_dout_12_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_inst_dout_13_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_inst_dout_13_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_inst_dout_14_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_inst_dout_14_rsci_iswt0
      = fsm_output[1];
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_inst_core_wten;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_inst_core_wten
      = ~ core_wen;
  wire [0:0] nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_inst_dout_15_rsci_iswt0;
  assign nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_inst_dout_15_rsci_iswt0
      = fsm_output[1];
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(din_rsc_z),
      .din_rsc_vz(din_rsc_vz),
      .din_rsc_lz(din_rsc_lz),
      .core_wen(core_wen),
      .din_rsci_oswt(reg_din_rsci_ld_core_psct_cse),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_d_mxwt(din_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_inst
      (
      .dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_inst_core_wten[0:0]),
      .dout_0_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsci_1_inst_dout_0_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_inst
      (
      .dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_inst_core_wten[0:0]),
      .dout_1_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsci_1_inst_dout_1_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_inst
      (
      .dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_inst_core_wten[0:0]),
      .dout_2_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsci_1_inst_dout_2_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_inst
      (
      .dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_inst_core_wten[0:0]),
      .dout_3_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsci_1_inst_dout_3_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_inst
      (
      .dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_inst_core_wten[0:0]),
      .dout_4_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsci_1_inst_dout_4_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_inst
      (
      .dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_inst_core_wten[0:0]),
      .dout_5_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsci_1_inst_dout_5_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_inst
      (
      .dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_inst_core_wten[0:0]),
      .dout_6_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsci_1_inst_dout_6_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_inst
      (
      .dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_inst_core_wten[0:0]),
      .dout_7_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsci_1_inst_dout_7_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_inst
      (
      .dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_inst_core_wten[0:0]),
      .dout_8_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsci_1_inst_dout_8_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_inst
      (
      .dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_inst_core_wten[0:0]),
      .dout_9_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsci_1_inst_dout_9_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_inst
      (
      .dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_inst_core_wten[0:0]),
      .dout_10_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsci_1_inst_dout_10_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_inst
      (
      .dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_inst_core_wten[0:0]),
      .dout_11_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsci_1_inst_dout_11_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_inst
      (
      .dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_inst_core_wten[0:0]),
      .dout_12_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsci_1_inst_dout_12_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_inst
      (
      .dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_inst_core_wten[0:0]),
      .dout_13_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsci_1_inst_dout_13_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_inst
      (
      .dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_inst_core_wten[0:0]),
      .dout_14_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsci_1_inst_dout_14_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_inst
      (
      .dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .core_wten(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_inst_core_wten[0:0]),
      .dout_15_rsci_iswt0(nl_WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsci_1_inst_dout_15_rsci_iswt0[0:0])
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_rls_obj_inst
      (
      .dout_15_rsc_rls_lz(dout_15_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_15_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_rls_obj_inst
      (
      .dout_14_rsc_rls_lz(dout_14_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_14_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_rls_obj_inst
      (
      .dout_13_rsc_rls_lz(dout_13_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_13_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_rls_obj_inst
      (
      .dout_12_rsc_rls_lz(dout_12_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_12_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_rls_obj_inst
      (
      .dout_11_rsc_rls_lz(dout_11_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_11_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_rls_obj_inst
      (
      .dout_10_rsc_rls_lz(dout_10_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_10_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_rls_obj_inst
      (
      .dout_9_rsc_rls_lz(dout_9_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_9_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_rls_obj_inst
      (
      .dout_8_rsc_rls_lz(dout_8_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_8_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_rls_obj_inst
      (
      .dout_7_rsc_rls_lz(dout_7_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_7_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_rls_obj_inst
      (
      .dout_6_rsc_rls_lz(dout_6_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_6_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_rls_obj_inst
      (
      .dout_5_rsc_rls_lz(dout_5_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_5_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_rls_obj_inst
      (
      .dout_4_rsc_rls_lz(dout_4_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_4_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_rls_obj_inst
      (
      .dout_3_rsc_rls_lz(dout_3_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_3_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_rls_obj_inst
      (
      .dout_2_rsc_rls_lz(dout_2_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_2_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_rls_obj_inst
      (
      .dout_1_rsc_rls_lz(dout_1_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_1_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_rls_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_rls_obj_inst
      (
      .dout_0_rsc_rls_lz(dout_0_rsc_rls_lz),
      .core_wten(core_wten),
      .dout_0_rsc_rls_obj_iswt0(reg_dout_0_rsc_rls_obj_ld_core_psct_cse)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_15_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_15_rsc_req_vz(dout_15_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_15_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_15_rsc_req_obj_wen_comp(dout_15_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_14_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_14_rsc_req_vz(dout_14_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_14_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_14_rsc_req_obj_wen_comp(dout_14_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_13_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_13_rsc_req_vz(dout_13_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_13_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_13_rsc_req_obj_wen_comp(dout_13_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_12_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_12_rsc_req_vz(dout_12_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_12_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_12_rsc_req_obj_wen_comp(dout_12_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_11_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_11_rsc_req_vz(dout_11_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_11_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_11_rsc_req_obj_wen_comp(dout_11_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_10_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_10_rsc_req_vz(dout_10_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_10_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_10_rsc_req_obj_wen_comp(dout_10_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_9_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_9_rsc_req_vz(dout_9_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_9_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_9_rsc_req_obj_wen_comp(dout_9_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_8_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_8_rsc_req_vz(dout_8_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_8_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_8_rsc_req_obj_wen_comp(dout_8_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_7_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_7_rsc_req_vz(dout_7_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_7_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_7_rsc_req_obj_wen_comp(dout_7_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_6_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_6_rsc_req_vz(dout_6_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_6_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_6_rsc_req_obj_wen_comp(dout_6_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_5_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_5_rsc_req_vz(dout_5_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_5_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_5_rsc_req_obj_wen_comp(dout_5_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_4_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_4_rsc_req_vz(dout_4_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_4_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_4_rsc_req_obj_wen_comp(dout_4_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_3_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_3_rsc_req_vz(dout_3_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_3_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_3_rsc_req_obj_wen_comp(dout_3_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_2_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_2_rsc_req_vz(dout_2_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_2_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_2_rsc_req_obj_wen_comp(dout_2_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_1_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_1_rsc_req_vz(dout_1_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_1_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_1_rsc_req_obj_wen_comp(dout_1_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_0_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_0_rsc_req_vz(dout_0_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_0_rsc_req_obj_oswt(reg_dout_15_rsc_req_obj_oswt_cse),
      .dout_0_rsc_req_obj_wen_comp(dout_0_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_staller WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .core_wten(core_wten),
      .dout_15_rsc_req_obj_wen_comp(dout_15_rsc_req_obj_wen_comp),
      .dout_14_rsc_req_obj_wen_comp(dout_14_rsc_req_obj_wen_comp),
      .dout_13_rsc_req_obj_wen_comp(dout_13_rsc_req_obj_wen_comp),
      .dout_12_rsc_req_obj_wen_comp(dout_12_rsc_req_obj_wen_comp),
      .dout_11_rsc_req_obj_wen_comp(dout_11_rsc_req_obj_wen_comp),
      .dout_10_rsc_req_obj_wen_comp(dout_10_rsc_req_obj_wen_comp),
      .dout_9_rsc_req_obj_wen_comp(dout_9_rsc_req_obj_wen_comp),
      .dout_8_rsc_req_obj_wen_comp(dout_8_rsc_req_obj_wen_comp),
      .dout_7_rsc_req_obj_wen_comp(dout_7_rsc_req_obj_wen_comp),
      .dout_6_rsc_req_obj_wen_comp(dout_6_rsc_req_obj_wen_comp),
      .dout_5_rsc_req_obj_wen_comp(dout_5_rsc_req_obj_wen_comp),
      .dout_4_rsc_req_obj_wen_comp(dout_4_rsc_req_obj_wen_comp),
      .dout_3_rsc_req_obj_wen_comp(dout_3_rsc_req_obj_wen_comp),
      .dout_2_rsc_req_obj_wen_comp(dout_2_rsc_req_obj_wen_comp),
      .dout_1_rsc_req_obj_wen_comp(dout_1_rsc_req_obj_wen_comp),
      .dout_0_rsc_req_obj_wen_comp(dout_0_rsc_req_obj_wen_comp)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign for_and_cse = core_wen & (~ (fsm_output[0]));
  assign WRITE_y_idx_and_cse = core_wen & nand_1_cse;
  assign nand_1_cse = ~((WRITE_acc_17_tmp[6]) & (for_k_idx_2_0_sva_1[2]));
  assign nor_nl = ~(exit_for_lpi_1_dfm_2 | exitL_exit_for_sva);
  assign WRITE_y_idx_6_0_lpi_1_dfm_5_0 = MUX_v_6_2_2(6'b000000, WRITE_y_idx_6_0_lpi_1_dfm_2_5_0_2,
      (nor_nl));
  assign for_not_7_nl = ~ exitL_exit_for_sva;
  assign for_k_idx_2_0_lpi_1_dfm_1_0 = MUX_v_2_2_2(2'b00, for_k_idx_2_0_lpi_1_dfm_1_1_0_1,
      (for_not_7_nl));
  assign exit_for_lpi_1_dfm_2_mx0w0 = (for_k_idx_2_0_sva_1[2]) & (WRITE_acc_17_tmp[6]);
  assign nl_for_k_idx_2_0_sva_1 = conv_u2u_2_3(for_k_idx_2_0_lpi_1_dfm_1_0) + 3'b1;
  assign for_k_idx_2_0_sva_1 = nl_for_k_idx_2_0_sva_1[2:0];
  assign nl_WRITE_acc_17_tmp = conv_u2u_6_7(WRITE_y_idx_6_0_lpi_1_dfm_5_0) + 7'b1;
  assign WRITE_acc_17_tmp = nl_WRITE_acc_17_tmp[6:0];
  assign dout_0_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_0_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_0_rsci_dinb_d = din_rsci_d_mxwt[63:0];
  assign dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_1_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_1_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_1_rsci_dinb_d = din_rsci_d_mxwt[127:64];
  assign dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_2_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_2_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_2_rsci_dinb_d = din_rsci_d_mxwt[191:128];
  assign dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_3_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_3_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_3_rsci_dinb_d = din_rsci_d_mxwt[255:192];
  assign dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_4_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_4_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_4_rsci_dinb_d = din_rsci_d_mxwt[319:256];
  assign dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_5_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_5_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_5_rsci_dinb_d = din_rsci_d_mxwt[383:320];
  assign dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_6_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_6_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_6_rsci_dinb_d = din_rsci_d_mxwt[447:384];
  assign dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_7_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_7_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_7_rsci_dinb_d = din_rsci_d_mxwt[511:448];
  assign dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_8_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_8_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_8_rsci_dinb_d = din_rsci_d_mxwt[575:512];
  assign dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_9_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_9_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_9_rsci_dinb_d = din_rsci_d_mxwt[639:576];
  assign dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_10_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_10_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_10_rsci_dinb_d = din_rsci_d_mxwt[703:640];
  assign dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_11_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_11_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_11_rsci_dinb_d = din_rsci_d_mxwt[767:704];
  assign dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_12_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_12_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_12_rsci_dinb_d = din_rsci_d_mxwt[831:768];
  assign dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_13_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_13_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_13_rsci_dinb_d = din_rsci_d_mxwt[895:832];
  assign dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_14_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_14_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_14_rsci_dinb_d = din_rsci_d_mxwt[959:896];
  assign dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign dout_15_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_15_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , WRITE_y_idx_6_0_lpi_1_dfm_5_0};
  assign dout_15_rsci_dinb_d = din_rsci_d_mxwt[1023:960];
  assign dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      reg_dout_15_rsc_req_obj_oswt_cse <= 1'b0;
      reg_dout_0_rsc_rls_obj_ld_core_psct_cse <= 1'b0;
      reg_din_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_dout_15_rsc_req_obj_oswt_cse <= ~(nand_1_cse & (fsm_output[1]));
      reg_dout_0_rsc_rls_obj_ld_core_psct_cse <= (WRITE_acc_17_tmp[6]) & (for_k_idx_2_0_sva_1[2])
          & (fsm_output[1]);
      reg_din_rsci_ld_core_psct_cse <= 1'b1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exitL_exit_for_sva <= 1'b1;
      exit_for_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( for_and_cse ) begin
      exitL_exit_for_sva <= exit_for_lpi_1_dfm_2_mx0w0;
      exit_for_lpi_1_dfm_2 <= exit_for_lpi_1_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      WRITE_y_idx_6_0_lpi_1_dfm_2_5_0_2 <= 6'b0;
      for_k_idx_2_0_lpi_1_dfm_1_1_0_1 <= 2'b0;
    end
    else if ( WRITE_y_idx_and_cse ) begin
      WRITE_y_idx_6_0_lpi_1_dfm_2_5_0_2 <= WRITE_acc_17_tmp[5:0];
      for_k_idx_2_0_lpi_1_dfm_1_1_0_1 <= MUX_v_2_2_2(for_k_idx_2_0_lpi_1_dfm_1_0,
          (for_k_idx_2_0_sva_1[1:0]), WRITE_acc_17_tmp[6]);
    end
  end

  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function  [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core (
  clk, rst, din_0_rsc_req_vz, din_0_rsc_rls_lz, din_1_rsc_req_vz, din_1_rsc_rls_lz,
      din_2_rsc_req_vz, din_2_rsc_rls_lz, din_3_rsc_req_vz, din_3_rsc_rls_lz, din_4_rsc_req_vz,
      din_4_rsc_rls_lz, din_5_rsc_req_vz, din_5_rsc_rls_lz, din_6_rsc_req_vz, din_6_rsc_rls_lz,
      din_7_rsc_req_vz, din_7_rsc_rls_lz, din_8_rsc_req_vz, din_8_rsc_rls_lz, din_9_rsc_req_vz,
      din_9_rsc_rls_lz, din_10_rsc_req_vz, din_10_rsc_rls_lz, din_11_rsc_req_vz,
      din_11_rsc_rls_lz, din_12_rsc_req_vz, din_12_rsc_rls_lz, din_13_rsc_req_vz,
      din_13_rsc_rls_lz, din_14_rsc_req_vz, din_14_rsc_rls_lz, din_15_rsc_req_vz,
      din_15_rsc_rls_lz, dout_rsc_z, dout_rsc_vz, dout_rsc_lz, din_0_rsci_addra_d,
      din_0_rsci_addrb_d, din_0_rsci_douta_d, din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_1_rsci_addra_d, din_1_rsci_addrb_d, din_1_rsci_douta_d, din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_2_rsci_addra_d, din_2_rsci_addrb_d, din_2_rsci_douta_d, din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_3_rsci_addra_d, din_3_rsci_addrb_d, din_3_rsci_douta_d, din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_4_rsci_addra_d, din_4_rsci_addrb_d, din_4_rsci_douta_d, din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_5_rsci_addra_d, din_5_rsci_addrb_d, din_5_rsci_douta_d, din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_6_rsci_addra_d, din_6_rsci_addrb_d, din_6_rsci_douta_d, din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_7_rsci_addra_d, din_7_rsci_addrb_d, din_7_rsci_douta_d, din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_8_rsci_addra_d, din_8_rsci_addrb_d, din_8_rsci_douta_d, din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_9_rsci_addra_d, din_9_rsci_addrb_d, din_9_rsci_douta_d, din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_10_rsci_addra_d, din_10_rsci_addrb_d, din_10_rsci_douta_d, din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_11_rsci_addra_d, din_11_rsci_addrb_d, din_11_rsci_douta_d, din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_12_rsci_addra_d, din_12_rsci_addrb_d, din_12_rsci_douta_d, din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_13_rsci_addra_d, din_13_rsci_addrb_d, din_13_rsci_douta_d, din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_14_rsci_addra_d, din_14_rsci_addrb_d, din_14_rsci_douta_d, din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      din_15_rsci_addra_d, din_15_rsci_addrb_d, din_15_rsci_douta_d, din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d
);
  input clk;
  input rst;
  input din_0_rsc_req_vz;
  output din_0_rsc_rls_lz;
  input din_1_rsc_req_vz;
  output din_1_rsc_rls_lz;
  input din_2_rsc_req_vz;
  output din_2_rsc_rls_lz;
  input din_3_rsc_req_vz;
  output din_3_rsc_rls_lz;
  input din_4_rsc_req_vz;
  output din_4_rsc_rls_lz;
  input din_5_rsc_req_vz;
  output din_5_rsc_rls_lz;
  input din_6_rsc_req_vz;
  output din_6_rsc_rls_lz;
  input din_7_rsc_req_vz;
  output din_7_rsc_rls_lz;
  input din_8_rsc_req_vz;
  output din_8_rsc_rls_lz;
  input din_9_rsc_req_vz;
  output din_9_rsc_rls_lz;
  input din_10_rsc_req_vz;
  output din_10_rsc_rls_lz;
  input din_11_rsc_req_vz;
  output din_11_rsc_rls_lz;
  input din_12_rsc_req_vz;
  output din_12_rsc_rls_lz;
  input din_13_rsc_req_vz;
  output din_13_rsc_rls_lz;
  input din_14_rsc_req_vz;
  output din_14_rsc_rls_lz;
  input din_15_rsc_req_vz;
  output din_15_rsc_rls_lz;
  output [1023:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;
  output [7:0] din_0_rsci_addra_d;
  output [7:0] din_0_rsci_addrb_d;
  input [63:0] din_0_rsci_douta_d;
  output din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_1_rsci_addra_d;
  output [7:0] din_1_rsci_addrb_d;
  input [63:0] din_1_rsci_douta_d;
  output din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_2_rsci_addra_d;
  output [7:0] din_2_rsci_addrb_d;
  input [63:0] din_2_rsci_douta_d;
  output din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_3_rsci_addra_d;
  output [7:0] din_3_rsci_addrb_d;
  input [63:0] din_3_rsci_douta_d;
  output din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_4_rsci_addra_d;
  output [7:0] din_4_rsci_addrb_d;
  input [63:0] din_4_rsci_douta_d;
  output din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_5_rsci_addra_d;
  output [7:0] din_5_rsci_addrb_d;
  input [63:0] din_5_rsci_douta_d;
  output din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_6_rsci_addra_d;
  output [7:0] din_6_rsci_addrb_d;
  input [63:0] din_6_rsci_douta_d;
  output din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_7_rsci_addra_d;
  output [7:0] din_7_rsci_addrb_d;
  input [63:0] din_7_rsci_douta_d;
  output din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_8_rsci_addra_d;
  output [7:0] din_8_rsci_addrb_d;
  input [63:0] din_8_rsci_douta_d;
  output din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_9_rsci_addra_d;
  output [7:0] din_9_rsci_addrb_d;
  input [63:0] din_9_rsci_douta_d;
  output din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_10_rsci_addra_d;
  output [7:0] din_10_rsci_addrb_d;
  input [63:0] din_10_rsci_douta_d;
  output din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_11_rsci_addra_d;
  output [7:0] din_11_rsci_addrb_d;
  input [63:0] din_11_rsci_douta_d;
  output din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_12_rsci_addra_d;
  output [7:0] din_12_rsci_addrb_d;
  input [63:0] din_12_rsci_douta_d;
  output din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_13_rsci_addra_d;
  output [7:0] din_13_rsci_addrb_d;
  input [63:0] din_13_rsci_douta_d;
  output din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_14_rsci_addra_d;
  output [7:0] din_14_rsci_addrb_d;
  input [63:0] din_14_rsci_douta_d;
  output din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] din_15_rsci_addra_d;
  output [7:0] din_15_rsci_addrb_d;
  input [63:0] din_15_rsci_douta_d;
  output din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations
  wire core_wen;
  wire [63:0] din_0_rsci_douta_d_mxwt;
  wire core_wten;
  wire [63:0] din_1_rsci_douta_d_mxwt;
  wire [63:0] din_2_rsci_douta_d_mxwt;
  wire [63:0] din_3_rsci_douta_d_mxwt;
  wire [63:0] din_4_rsci_douta_d_mxwt;
  wire [63:0] din_5_rsci_douta_d_mxwt;
  wire [63:0] din_6_rsci_douta_d_mxwt;
  wire [63:0] din_7_rsci_douta_d_mxwt;
  wire [63:0] din_8_rsci_douta_d_mxwt;
  wire [63:0] din_9_rsci_douta_d_mxwt;
  wire [63:0] din_10_rsci_douta_d_mxwt;
  wire [63:0] din_11_rsci_douta_d_mxwt;
  wire [63:0] din_12_rsci_douta_d_mxwt;
  wire [63:0] din_13_rsci_douta_d_mxwt;
  wire [63:0] din_14_rsci_douta_d_mxwt;
  wire [63:0] din_15_rsci_douta_d_mxwt;
  wire dout_rsci_wen_comp;
  wire din_15_rsc_req_obj_wen_comp;
  wire din_14_rsc_req_obj_wen_comp;
  wire din_13_rsc_req_obj_wen_comp;
  wire din_12_rsc_req_obj_wen_comp;
  wire din_11_rsc_req_obj_wen_comp;
  wire din_10_rsc_req_obj_wen_comp;
  wire din_9_rsc_req_obj_wen_comp;
  wire din_8_rsc_req_obj_wen_comp;
  wire din_7_rsc_req_obj_wen_comp;
  wire din_6_rsc_req_obj_wen_comp;
  wire din_5_rsc_req_obj_wen_comp;
  wire din_4_rsc_req_obj_wen_comp;
  wire din_3_rsc_req_obj_wen_comp;
  wire din_2_rsc_req_obj_wen_comp;
  wire din_1_rsc_req_obj_wen_comp;
  wire din_0_rsc_req_obj_wen_comp;
  reg [63:0] dout_rsci_d_1023_960;
  reg [63:0] dout_rsci_d_959_896;
  reg [63:0] dout_rsci_d_895_832;
  reg [63:0] dout_rsci_d_831_768;
  reg [63:0] dout_rsci_d_767_704;
  reg [63:0] dout_rsci_d_703_640;
  reg [63:0] dout_rsci_d_639_576;
  reg [63:0] dout_rsci_d_575_512;
  reg [63:0] dout_rsci_d_511_448;
  reg [63:0] dout_rsci_d_447_384;
  reg [63:0] dout_rsci_d_383_320;
  reg [63:0] dout_rsci_d_319_256;
  reg [63:0] dout_rsci_d_255_192;
  reg [63:0] dout_rsci_d_191_128;
  reg [63:0] dout_rsci_d_127_64;
  reg [63:0] dout_rsci_d_63_0;
  wire [1:0] fsm_output;
  wire [6:0] READ_acc_33_tmp;
  wire [7:0] nl_READ_acc_33_tmp;
  reg exitL_exit_for_sva;
  reg exit_for_lpi_1_dfm_2;
  reg [1:0] for_k_idx_2_0_lpi_1_dfm_1_1_0_1;
  reg [5:0] READ_y_idx_6_0_lpi_1_dfm_2_5_0_2;
  wire [2:0] for_k_idx_2_0_sva_1;
  wire [3:0] nl_for_k_idx_2_0_sva_1;
  reg reg_din_15_rsc_req_obj_oswt_cse;
  wire dout_and_cse;
  reg reg_din_15_rsc_rls_obj_ld_core_psct_cse;
  reg reg_dout_rsci_ld_core_psct_cse;
  reg reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse;
  wire for_and_cse;
  wire nand_1_cse;
  wire din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire [1:0] for_k_idx_2_0_lpi_1_dfm_1_0;
  wire [5:0] READ_y_idx_6_0_lpi_1_dfm_5_0;
  wire exit_for_lpi_1_dfm_2_mx0w0;
  wire READ_y_idx_and_cse;

  wire[0:0] nor_nl;
  wire[0:0] for_not_7_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_inst_din_0_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_inst_din_0_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_inst_din_1_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_inst_din_1_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_inst_din_2_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_inst_din_2_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_inst_din_3_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_inst_din_3_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_inst_din_4_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_inst_din_4_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_inst_din_5_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_inst_din_5_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_inst_din_6_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_inst_din_6_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_inst_din_7_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_inst_din_7_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_inst_din_8_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_inst_din_8_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_inst_din_9_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_inst_din_9_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_inst_din_10_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_inst_din_10_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_inst_din_11_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_inst_din_11_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_inst_din_12_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_inst_din_12_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_inst_din_13_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_inst_din_13_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_inst_din_14_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_inst_din_14_rsci_oswt_pff
      = fsm_output[1];
  wire [0:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_inst_din_15_rsci_oswt_pff;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_inst_din_15_rsci_oswt_pff
      = fsm_output[1];
  wire [1023:0] nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_inst_dout_rsci_d;
  assign nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_inst_dout_rsci_d = {dout_rsci_d_1023_960
      , dout_rsci_d_959_896 , dout_rsci_d_895_832 , dout_rsci_d_831_768 , dout_rsci_d_767_704
      , dout_rsci_d_703_640 , dout_rsci_d_639_576 , dout_rsci_d_575_512 , dout_rsci_d_511_448
      , dout_rsci_d_447_384 , dout_rsci_d_383_320 , dout_rsci_d_319_256 , dout_rsci_d_255_192
      , dout_rsci_d_191_128 , dout_rsci_d_127_64 , dout_rsci_d_63_0};
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_0_rsci_douta_d(din_0_rsci_douta_d),
      .din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .din_0_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_0_rsci_douta_d_mxwt(din_0_rsci_douta_d_mxwt),
      .core_wten(core_wten),
      .din_0_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsci_1_inst_din_0_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_1_rsci_douta_d(din_1_rsci_douta_d),
      .din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_1_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_1_rsci_douta_d_mxwt(din_1_rsci_douta_d_mxwt),
      .din_1_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsci_1_inst_din_1_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_2_rsci_douta_d(din_2_rsci_douta_d),
      .din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_2_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_2_rsci_douta_d_mxwt(din_2_rsci_douta_d_mxwt),
      .din_2_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsci_1_inst_din_2_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_3_rsci_douta_d(din_3_rsci_douta_d),
      .din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_3_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_3_rsci_douta_d_mxwt(din_3_rsci_douta_d_mxwt),
      .din_3_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsci_1_inst_din_3_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_4_rsci_douta_d(din_4_rsci_douta_d),
      .din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_4_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_4_rsci_douta_d_mxwt(din_4_rsci_douta_d_mxwt),
      .din_4_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsci_1_inst_din_4_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_5_rsci_douta_d(din_5_rsci_douta_d),
      .din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_5_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_5_rsci_douta_d_mxwt(din_5_rsci_douta_d_mxwt),
      .din_5_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsci_1_inst_din_5_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_6_rsci_douta_d(din_6_rsci_douta_d),
      .din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_6_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_6_rsci_douta_d_mxwt(din_6_rsci_douta_d_mxwt),
      .din_6_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsci_1_inst_din_6_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_7_rsci_douta_d(din_7_rsci_douta_d),
      .din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_7_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_7_rsci_douta_d_mxwt(din_7_rsci_douta_d_mxwt),
      .din_7_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsci_1_inst_din_7_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_8_rsci_douta_d(din_8_rsci_douta_d),
      .din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_8_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_8_rsci_douta_d_mxwt(din_8_rsci_douta_d_mxwt),
      .din_8_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsci_1_inst_din_8_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_9_rsci_douta_d(din_9_rsci_douta_d),
      .din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_9_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_9_rsci_douta_d_mxwt(din_9_rsci_douta_d_mxwt),
      .din_9_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsci_1_inst_din_9_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_10_rsci_douta_d(din_10_rsci_douta_d),
      .din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_10_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_10_rsci_douta_d_mxwt(din_10_rsci_douta_d_mxwt),
      .din_10_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsci_1_inst_din_10_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_11_rsci_douta_d(din_11_rsci_douta_d),
      .din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_11_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_11_rsci_douta_d_mxwt(din_11_rsci_douta_d_mxwt),
      .din_11_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsci_1_inst_din_11_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_12_rsci_douta_d(din_12_rsci_douta_d),
      .din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_12_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_12_rsci_douta_d_mxwt(din_12_rsci_douta_d_mxwt),
      .din_12_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsci_1_inst_din_12_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_13_rsci_douta_d(din_13_rsci_douta_d),
      .din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_13_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_13_rsci_douta_d_mxwt(din_13_rsci_douta_d_mxwt),
      .din_13_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsci_1_inst_din_13_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_14_rsci_douta_d(din_14_rsci_douta_d),
      .din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_14_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_14_rsci_douta_d_mxwt(din_14_rsci_douta_d_mxwt),
      .din_14_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsci_1_inst_din_14_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .din_15_rsci_douta_d(din_15_rsci_douta_d),
      .din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_15_rsci_oswt(reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .din_15_rsci_douta_d_mxwt(din_15_rsci_douta_d_mxwt),
      .din_15_rsci_oswt_pff(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsci_1_inst_din_15_rsci_oswt_pff[0:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dout_rsc_z(dout_rsc_z),
      .dout_rsc_vz(dout_rsc_vz),
      .dout_rsc_lz(dout_rsc_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsci_oswt(reg_dout_rsci_ld_core_psct_cse),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_d(nl_READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_dout_rsci_inst_dout_rsci_d[1023:0])
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_rls_obj_inst
      (
      .din_0_rsc_rls_lz(din_0_rsc_rls_lz),
      .core_wten(core_wten),
      .din_0_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_rls_obj_inst
      (
      .din_1_rsc_rls_lz(din_1_rsc_rls_lz),
      .core_wten(core_wten),
      .din_1_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_rls_obj_inst
      (
      .din_2_rsc_rls_lz(din_2_rsc_rls_lz),
      .core_wten(core_wten),
      .din_2_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_rls_obj_inst
      (
      .din_3_rsc_rls_lz(din_3_rsc_rls_lz),
      .core_wten(core_wten),
      .din_3_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_rls_obj_inst
      (
      .din_4_rsc_rls_lz(din_4_rsc_rls_lz),
      .core_wten(core_wten),
      .din_4_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_rls_obj_inst
      (
      .din_5_rsc_rls_lz(din_5_rsc_rls_lz),
      .core_wten(core_wten),
      .din_5_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_rls_obj_inst
      (
      .din_6_rsc_rls_lz(din_6_rsc_rls_lz),
      .core_wten(core_wten),
      .din_6_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_rls_obj_inst
      (
      .din_7_rsc_rls_lz(din_7_rsc_rls_lz),
      .core_wten(core_wten),
      .din_7_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_rls_obj_inst
      (
      .din_8_rsc_rls_lz(din_8_rsc_rls_lz),
      .core_wten(core_wten),
      .din_8_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_rls_obj_inst
      (
      .din_9_rsc_rls_lz(din_9_rsc_rls_lz),
      .core_wten(core_wten),
      .din_9_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_rls_obj_inst
      (
      .din_10_rsc_rls_lz(din_10_rsc_rls_lz),
      .core_wten(core_wten),
      .din_10_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_rls_obj_inst
      (
      .din_11_rsc_rls_lz(din_11_rsc_rls_lz),
      .core_wten(core_wten),
      .din_11_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_rls_obj_inst
      (
      .din_12_rsc_rls_lz(din_12_rsc_rls_lz),
      .core_wten(core_wten),
      .din_12_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_rls_obj_inst
      (
      .din_13_rsc_rls_lz(din_13_rsc_rls_lz),
      .core_wten(core_wten),
      .din_13_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_rls_obj_inst
      (
      .din_14_rsc_rls_lz(din_14_rsc_rls_lz),
      .core_wten(core_wten),
      .din_14_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_rls_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_rls_obj_inst
      (
      .din_15_rsc_rls_lz(din_15_rsc_rls_lz),
      .core_wten(core_wten),
      .din_15_rsc_rls_obj_iswt0(reg_din_15_rsc_rls_obj_ld_core_psct_cse)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_15_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_15_rsc_req_vz(din_15_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_15_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_15_rsc_req_obj_wen_comp(din_15_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_14_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_14_rsc_req_vz(din_14_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_14_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_14_rsc_req_obj_wen_comp(din_14_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_13_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_13_rsc_req_vz(din_13_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_13_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_13_rsc_req_obj_wen_comp(din_13_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_12_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_12_rsc_req_vz(din_12_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_12_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_12_rsc_req_obj_wen_comp(din_12_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_11_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_11_rsc_req_vz(din_11_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_11_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_11_rsc_req_obj_wen_comp(din_11_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_10_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_10_rsc_req_vz(din_10_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_10_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_10_rsc_req_obj_wen_comp(din_10_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_9_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_9_rsc_req_vz(din_9_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_9_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_9_rsc_req_obj_wen_comp(din_9_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_8_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_8_rsc_req_vz(din_8_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_8_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_8_rsc_req_obj_wen_comp(din_8_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_7_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_7_rsc_req_vz(din_7_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_7_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_7_rsc_req_obj_wen_comp(din_7_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_6_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_6_rsc_req_vz(din_6_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_6_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_6_rsc_req_obj_wen_comp(din_6_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_5_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_5_rsc_req_vz(din_5_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_5_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_5_rsc_req_obj_wen_comp(din_5_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_4_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_4_rsc_req_vz(din_4_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_4_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_4_rsc_req_obj_wen_comp(din_4_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_3_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_3_rsc_req_vz(din_3_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_3_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_3_rsc_req_obj_wen_comp(din_3_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_2_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_2_rsc_req_vz(din_2_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_2_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_2_rsc_req_obj_wen_comp(din_2_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_1_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_1_rsc_req_vz(din_1_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_1_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_1_rsc_req_obj_wen_comp(din_1_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_din_0_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .din_0_rsc_req_vz(din_0_rsc_req_vz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .din_0_rsc_req_obj_oswt(reg_din_15_rsc_req_obj_oswt_cse),
      .din_0_rsc_req_obj_wen_comp(din_0_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_staller READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .din_15_rsc_req_obj_wen_comp(din_15_rsc_req_obj_wen_comp),
      .din_14_rsc_req_obj_wen_comp(din_14_rsc_req_obj_wen_comp),
      .din_13_rsc_req_obj_wen_comp(din_13_rsc_req_obj_wen_comp),
      .din_12_rsc_req_obj_wen_comp(din_12_rsc_req_obj_wen_comp),
      .din_11_rsc_req_obj_wen_comp(din_11_rsc_req_obj_wen_comp),
      .din_10_rsc_req_obj_wen_comp(din_10_rsc_req_obj_wen_comp),
      .din_9_rsc_req_obj_wen_comp(din_9_rsc_req_obj_wen_comp),
      .din_8_rsc_req_obj_wen_comp(din_8_rsc_req_obj_wen_comp),
      .din_7_rsc_req_obj_wen_comp(din_7_rsc_req_obj_wen_comp),
      .din_6_rsc_req_obj_wen_comp(din_6_rsc_req_obj_wen_comp),
      .din_5_rsc_req_obj_wen_comp(din_5_rsc_req_obj_wen_comp),
      .din_4_rsc_req_obj_wen_comp(din_4_rsc_req_obj_wen_comp),
      .din_3_rsc_req_obj_wen_comp(din_3_rsc_req_obj_wen_comp),
      .din_2_rsc_req_obj_wen_comp(din_2_rsc_req_obj_wen_comp),
      .din_1_rsc_req_obj_wen_comp(din_1_rsc_req_obj_wen_comp),
      .din_0_rsc_req_obj_wen_comp(din_0_rsc_req_obj_wen_comp)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_core_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign dout_and_cse = core_wen & reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse;
  assign for_and_cse = core_wen & (~ (fsm_output[0]));
  assign READ_y_idx_and_cse = core_wen & nand_1_cse;
  assign nand_1_cse = ~((READ_acc_33_tmp[6]) & (for_k_idx_2_0_sva_1[2]));
  assign nor_nl = ~(exit_for_lpi_1_dfm_2 | exitL_exit_for_sva);
  assign READ_y_idx_6_0_lpi_1_dfm_5_0 = MUX_v_6_2_2(6'b000000, READ_y_idx_6_0_lpi_1_dfm_2_5_0_2,
      (nor_nl));
  assign for_not_7_nl = ~ exitL_exit_for_sva;
  assign for_k_idx_2_0_lpi_1_dfm_1_0 = MUX_v_2_2_2(2'b00, for_k_idx_2_0_lpi_1_dfm_1_1_0_1,
      (for_not_7_nl));
  assign exit_for_lpi_1_dfm_2_mx0w0 = (for_k_idx_2_0_sva_1[2]) & (READ_acc_33_tmp[6]);
  assign nl_for_k_idx_2_0_sva_1 = conv_u2u_2_3(for_k_idx_2_0_lpi_1_dfm_1_0) + 3'b1;
  assign for_k_idx_2_0_sva_1 = nl_for_k_idx_2_0_sva_1[2:0];
  assign nl_READ_acc_33_tmp = conv_u2u_6_7(READ_y_idx_6_0_lpi_1_dfm_5_0) + 7'b1;
  assign READ_acc_33_tmp = nl_READ_acc_33_tmp[6:0];
  assign din_0_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_0_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_1_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_1_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_2_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_2_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_3_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_3_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_4_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_4_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_5_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_5_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_6_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_6_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_7_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_7_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_8_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_8_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_9_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_9_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_10_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_10_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_11_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_11_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_12_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_12_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_13_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_13_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_14_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_14_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign din_15_rsci_addra_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_15_rsci_addrb_d = {for_k_idx_2_0_lpi_1_dfm_1_0 , READ_y_idx_6_0_lpi_1_dfm_5_0};
  assign din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      reg_din_15_rsc_req_obj_oswt_cse <= 1'b0;
      reg_din_15_rsc_rls_obj_ld_core_psct_cse <= 1'b0;
      reg_dout_rsci_ld_core_psct_cse <= 1'b0;
      reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_din_15_rsc_req_obj_oswt_cse <= ~(nand_1_cse & (fsm_output[1]));
      reg_din_15_rsc_rls_obj_ld_core_psct_cse <= (READ_acc_33_tmp[6]) & (for_k_idx_2_0_sva_1[2])
          & (fsm_output[1]);
      reg_dout_rsci_ld_core_psct_cse <= reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse;
      reg_din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_core_psct_cse <= fsm_output[1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      dout_rsci_d_63_0 <= 64'b0;
      dout_rsci_d_127_64 <= 64'b0;
      dout_rsci_d_191_128 <= 64'b0;
      dout_rsci_d_255_192 <= 64'b0;
      dout_rsci_d_319_256 <= 64'b0;
      dout_rsci_d_383_320 <= 64'b0;
      dout_rsci_d_447_384 <= 64'b0;
      dout_rsci_d_511_448 <= 64'b0;
      dout_rsci_d_575_512 <= 64'b0;
      dout_rsci_d_639_576 <= 64'b0;
      dout_rsci_d_703_640 <= 64'b0;
      dout_rsci_d_767_704 <= 64'b0;
      dout_rsci_d_831_768 <= 64'b0;
      dout_rsci_d_895_832 <= 64'b0;
      dout_rsci_d_959_896 <= 64'b0;
      dout_rsci_d_1023_960 <= 64'b0;
    end
    else if ( dout_and_cse ) begin
      dout_rsci_d_63_0 <= din_0_rsci_douta_d_mxwt;
      dout_rsci_d_127_64 <= din_1_rsci_douta_d_mxwt;
      dout_rsci_d_191_128 <= din_2_rsci_douta_d_mxwt;
      dout_rsci_d_255_192 <= din_3_rsci_douta_d_mxwt;
      dout_rsci_d_319_256 <= din_4_rsci_douta_d_mxwt;
      dout_rsci_d_383_320 <= din_5_rsci_douta_d_mxwt;
      dout_rsci_d_447_384 <= din_6_rsci_douta_d_mxwt;
      dout_rsci_d_511_448 <= din_7_rsci_douta_d_mxwt;
      dout_rsci_d_575_512 <= din_8_rsci_douta_d_mxwt;
      dout_rsci_d_639_576 <= din_9_rsci_douta_d_mxwt;
      dout_rsci_d_703_640 <= din_10_rsci_douta_d_mxwt;
      dout_rsci_d_767_704 <= din_11_rsci_douta_d_mxwt;
      dout_rsci_d_831_768 <= din_12_rsci_douta_d_mxwt;
      dout_rsci_d_895_832 <= din_13_rsci_douta_d_mxwt;
      dout_rsci_d_959_896 <= din_14_rsci_douta_d_mxwt;
      dout_rsci_d_1023_960 <= din_15_rsci_douta_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exitL_exit_for_sva <= 1'b1;
      exit_for_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( for_and_cse ) begin
      exitL_exit_for_sva <= exit_for_lpi_1_dfm_2_mx0w0;
      exit_for_lpi_1_dfm_2 <= exit_for_lpi_1_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      READ_y_idx_6_0_lpi_1_dfm_2_5_0_2 <= 6'b0;
      for_k_idx_2_0_lpi_1_dfm_1_1_0_1 <= 2'b0;
    end
    else if ( READ_y_idx_and_cse ) begin
      READ_y_idx_6_0_lpi_1_dfm_2_5_0_2 <= READ_acc_33_tmp[5:0];
      for_k_idx_2_0_lpi_1_dfm_1_1_0_1 <= MUX_v_2_2_2(for_k_idx_2_0_lpi_1_dfm_1_0,
          (for_k_idx_2_0_sva_1[1:0]), READ_acc_33_tmp[6]);
    end
  end

  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function  [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_1
// ------------------------------------------------------------------


module WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_1 (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, dout_0_rsc_csa_n, dout_0_rsc_csb_n,
      dout_0_rsc_addra, dout_0_rsc_addrb, dout_0_rsc_dinb, dout_0_rsc_douta, dout_0_rsc_req_vz,
      dout_0_rsc_rls_lz, dout_1_rsc_csa_n, dout_1_rsc_csb_n, dout_1_rsc_addra, dout_1_rsc_addrb,
      dout_1_rsc_dinb, dout_1_rsc_douta, dout_1_rsc_req_vz, dout_1_rsc_rls_lz, dout_2_rsc_csa_n,
      dout_2_rsc_csb_n, dout_2_rsc_addra, dout_2_rsc_addrb, dout_2_rsc_dinb, dout_2_rsc_douta,
      dout_2_rsc_req_vz, dout_2_rsc_rls_lz, dout_3_rsc_csa_n, dout_3_rsc_csb_n, dout_3_rsc_addra,
      dout_3_rsc_addrb, dout_3_rsc_dinb, dout_3_rsc_douta, dout_3_rsc_req_vz, dout_3_rsc_rls_lz,
      dout_4_rsc_csa_n, dout_4_rsc_csb_n, dout_4_rsc_addra, dout_4_rsc_addrb, dout_4_rsc_dinb,
      dout_4_rsc_douta, dout_4_rsc_req_vz, dout_4_rsc_rls_lz, dout_5_rsc_csa_n, dout_5_rsc_csb_n,
      dout_5_rsc_addra, dout_5_rsc_addrb, dout_5_rsc_dinb, dout_5_rsc_douta, dout_5_rsc_req_vz,
      dout_5_rsc_rls_lz, dout_6_rsc_csa_n, dout_6_rsc_csb_n, dout_6_rsc_addra, dout_6_rsc_addrb,
      dout_6_rsc_dinb, dout_6_rsc_douta, dout_6_rsc_req_vz, dout_6_rsc_rls_lz, dout_7_rsc_csa_n,
      dout_7_rsc_csb_n, dout_7_rsc_addra, dout_7_rsc_addrb, dout_7_rsc_dinb, dout_7_rsc_douta,
      dout_7_rsc_req_vz, dout_7_rsc_rls_lz, dout_8_rsc_csa_n, dout_8_rsc_csb_n, dout_8_rsc_addra,
      dout_8_rsc_addrb, dout_8_rsc_dinb, dout_8_rsc_douta, dout_8_rsc_req_vz, dout_8_rsc_rls_lz,
      dout_9_rsc_csa_n, dout_9_rsc_csb_n, dout_9_rsc_addra, dout_9_rsc_addrb, dout_9_rsc_dinb,
      dout_9_rsc_douta, dout_9_rsc_req_vz, dout_9_rsc_rls_lz, dout_10_rsc_csa_n,
      dout_10_rsc_csb_n, dout_10_rsc_addra, dout_10_rsc_addrb, dout_10_rsc_dinb,
      dout_10_rsc_douta, dout_10_rsc_req_vz, dout_10_rsc_rls_lz, dout_11_rsc_csa_n,
      dout_11_rsc_csb_n, dout_11_rsc_addra, dout_11_rsc_addrb, dout_11_rsc_dinb,
      dout_11_rsc_douta, dout_11_rsc_req_vz, dout_11_rsc_rls_lz, dout_12_rsc_csa_n,
      dout_12_rsc_csb_n, dout_12_rsc_addra, dout_12_rsc_addrb, dout_12_rsc_dinb,
      dout_12_rsc_douta, dout_12_rsc_req_vz, dout_12_rsc_rls_lz, dout_13_rsc_csa_n,
      dout_13_rsc_csb_n, dout_13_rsc_addra, dout_13_rsc_addrb, dout_13_rsc_dinb,
      dout_13_rsc_douta, dout_13_rsc_req_vz, dout_13_rsc_rls_lz, dout_14_rsc_csa_n,
      dout_14_rsc_csb_n, dout_14_rsc_addra, dout_14_rsc_addrb, dout_14_rsc_dinb,
      dout_14_rsc_douta, dout_14_rsc_req_vz, dout_14_rsc_rls_lz, dout_15_rsc_csa_n,
      dout_15_rsc_csb_n, dout_15_rsc_addra, dout_15_rsc_addrb, dout_15_rsc_dinb,
      dout_15_rsc_douta, dout_15_rsc_req_vz, dout_15_rsc_rls_lz, dout_16_rsc_csa_n,
      dout_16_rsc_csb_n, dout_16_rsc_addra, dout_16_rsc_addrb, dout_16_rsc_dinb,
      dout_16_rsc_douta, dout_16_rsc_req_vz, dout_16_rsc_rls_lz, dout_17_rsc_csa_n,
      dout_17_rsc_csb_n, dout_17_rsc_addra, dout_17_rsc_addrb, dout_17_rsc_dinb,
      dout_17_rsc_douta, dout_17_rsc_req_vz, dout_17_rsc_rls_lz, clamp_mem, scan_n,
      shift_n, slp_nret_n, slp_ret_n
);
  input clk;
  input rst;
  input [15:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  output dout_0_rsc_csa_n;
  output dout_0_rsc_csb_n;
  output [6:0] dout_0_rsc_addra;
  output [6:0] dout_0_rsc_addrb;
  output [63:0] dout_0_rsc_dinb;
  input [63:0] dout_0_rsc_douta;
  input dout_0_rsc_req_vz;
  output dout_0_rsc_rls_lz;
  output dout_1_rsc_csa_n;
  output dout_1_rsc_csb_n;
  output [6:0] dout_1_rsc_addra;
  output [6:0] dout_1_rsc_addrb;
  output [63:0] dout_1_rsc_dinb;
  input [63:0] dout_1_rsc_douta;
  input dout_1_rsc_req_vz;
  output dout_1_rsc_rls_lz;
  output dout_2_rsc_csa_n;
  output dout_2_rsc_csb_n;
  output [6:0] dout_2_rsc_addra;
  output [6:0] dout_2_rsc_addrb;
  output [63:0] dout_2_rsc_dinb;
  input [63:0] dout_2_rsc_douta;
  input dout_2_rsc_req_vz;
  output dout_2_rsc_rls_lz;
  output dout_3_rsc_csa_n;
  output dout_3_rsc_csb_n;
  output [6:0] dout_3_rsc_addra;
  output [6:0] dout_3_rsc_addrb;
  output [63:0] dout_3_rsc_dinb;
  input [63:0] dout_3_rsc_douta;
  input dout_3_rsc_req_vz;
  output dout_3_rsc_rls_lz;
  output dout_4_rsc_csa_n;
  output dout_4_rsc_csb_n;
  output [6:0] dout_4_rsc_addra;
  output [6:0] dout_4_rsc_addrb;
  output [63:0] dout_4_rsc_dinb;
  input [63:0] dout_4_rsc_douta;
  input dout_4_rsc_req_vz;
  output dout_4_rsc_rls_lz;
  output dout_5_rsc_csa_n;
  output dout_5_rsc_csb_n;
  output [6:0] dout_5_rsc_addra;
  output [6:0] dout_5_rsc_addrb;
  output [63:0] dout_5_rsc_dinb;
  input [63:0] dout_5_rsc_douta;
  input dout_5_rsc_req_vz;
  output dout_5_rsc_rls_lz;
  output dout_6_rsc_csa_n;
  output dout_6_rsc_csb_n;
  output [6:0] dout_6_rsc_addra;
  output [6:0] dout_6_rsc_addrb;
  output [63:0] dout_6_rsc_dinb;
  input [63:0] dout_6_rsc_douta;
  input dout_6_rsc_req_vz;
  output dout_6_rsc_rls_lz;
  output dout_7_rsc_csa_n;
  output dout_7_rsc_csb_n;
  output [6:0] dout_7_rsc_addra;
  output [6:0] dout_7_rsc_addrb;
  output [63:0] dout_7_rsc_dinb;
  input [63:0] dout_7_rsc_douta;
  input dout_7_rsc_req_vz;
  output dout_7_rsc_rls_lz;
  output dout_8_rsc_csa_n;
  output dout_8_rsc_csb_n;
  output [6:0] dout_8_rsc_addra;
  output [6:0] dout_8_rsc_addrb;
  output [63:0] dout_8_rsc_dinb;
  input [63:0] dout_8_rsc_douta;
  input dout_8_rsc_req_vz;
  output dout_8_rsc_rls_lz;
  output dout_9_rsc_csa_n;
  output dout_9_rsc_csb_n;
  output [6:0] dout_9_rsc_addra;
  output [6:0] dout_9_rsc_addrb;
  output [63:0] dout_9_rsc_dinb;
  input [63:0] dout_9_rsc_douta;
  input dout_9_rsc_req_vz;
  output dout_9_rsc_rls_lz;
  output dout_10_rsc_csa_n;
  output dout_10_rsc_csb_n;
  output [6:0] dout_10_rsc_addra;
  output [6:0] dout_10_rsc_addrb;
  output [63:0] dout_10_rsc_dinb;
  input [63:0] dout_10_rsc_douta;
  input dout_10_rsc_req_vz;
  output dout_10_rsc_rls_lz;
  output dout_11_rsc_csa_n;
  output dout_11_rsc_csb_n;
  output [6:0] dout_11_rsc_addra;
  output [6:0] dout_11_rsc_addrb;
  output [63:0] dout_11_rsc_dinb;
  input [63:0] dout_11_rsc_douta;
  input dout_11_rsc_req_vz;
  output dout_11_rsc_rls_lz;
  output dout_12_rsc_csa_n;
  output dout_12_rsc_csb_n;
  output [6:0] dout_12_rsc_addra;
  output [6:0] dout_12_rsc_addrb;
  output [63:0] dout_12_rsc_dinb;
  input [63:0] dout_12_rsc_douta;
  input dout_12_rsc_req_vz;
  output dout_12_rsc_rls_lz;
  output dout_13_rsc_csa_n;
  output dout_13_rsc_csb_n;
  output [6:0] dout_13_rsc_addra;
  output [6:0] dout_13_rsc_addrb;
  output [63:0] dout_13_rsc_dinb;
  input [63:0] dout_13_rsc_douta;
  input dout_13_rsc_req_vz;
  output dout_13_rsc_rls_lz;
  output dout_14_rsc_csa_n;
  output dout_14_rsc_csb_n;
  output [6:0] dout_14_rsc_addra;
  output [6:0] dout_14_rsc_addrb;
  output [63:0] dout_14_rsc_dinb;
  input [63:0] dout_14_rsc_douta;
  input dout_14_rsc_req_vz;
  output dout_14_rsc_rls_lz;
  output dout_15_rsc_csa_n;
  output dout_15_rsc_csb_n;
  output [6:0] dout_15_rsc_addra;
  output [6:0] dout_15_rsc_addrb;
  output [63:0] dout_15_rsc_dinb;
  input [63:0] dout_15_rsc_douta;
  input dout_15_rsc_req_vz;
  output dout_15_rsc_rls_lz;
  output dout_16_rsc_csa_n;
  output dout_16_rsc_csb_n;
  output [6:0] dout_16_rsc_addra;
  output [6:0] dout_16_rsc_addrb;
  output [63:0] dout_16_rsc_dinb;
  input [63:0] dout_16_rsc_douta;
  input dout_16_rsc_req_vz;
  output dout_16_rsc_rls_lz;
  output dout_17_rsc_csa_n;
  output dout_17_rsc_csb_n;
  output [6:0] dout_17_rsc_addra;
  output [6:0] dout_17_rsc_addrb;
  output [63:0] dout_17_rsc_dinb;
  input [63:0] dout_17_rsc_douta;
  input dout_17_rsc_req_vz;
  output dout_17_rsc_rls_lz;
  input clamp_mem;
  input scan_n;
  input shift_n;
  input slp_nret_n;
  input slp_ret_n;


  // Interconnect Declarations
  wire [63:0] dout_0_rsci_dinb_d;
  wire [63:0] dout_0_rsci_douta_d;
  wire dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_1_rsci_dinb_d;
  wire [63:0] dout_1_rsci_douta_d;
  wire dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_2_rsci_dinb_d;
  wire [63:0] dout_2_rsci_douta_d;
  wire dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_3_rsci_dinb_d;
  wire [63:0] dout_3_rsci_douta_d;
  wire dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_4_rsci_dinb_d;
  wire [63:0] dout_4_rsci_douta_d;
  wire dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_5_rsci_dinb_d;
  wire [63:0] dout_5_rsci_douta_d;
  wire dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_6_rsci_dinb_d;
  wire [63:0] dout_6_rsci_douta_d;
  wire dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_7_rsci_dinb_d;
  wire [63:0] dout_7_rsci_douta_d;
  wire dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_8_rsci_dinb_d;
  wire [63:0] dout_8_rsci_douta_d;
  wire dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_9_rsci_dinb_d;
  wire [63:0] dout_9_rsci_douta_d;
  wire dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_10_rsci_dinb_d;
  wire [63:0] dout_10_rsci_douta_d;
  wire dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_11_rsci_dinb_d;
  wire [63:0] dout_11_rsci_douta_d;
  wire dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_12_rsci_dinb_d;
  wire [63:0] dout_12_rsci_douta_d;
  wire dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_13_rsci_dinb_d;
  wire [63:0] dout_13_rsci_douta_d;
  wire dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_14_rsci_dinb_d;
  wire [63:0] dout_14_rsci_douta_d;
  wire dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_15_rsci_dinb_d;
  wire [63:0] dout_15_rsci_douta_d;
  wire dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_16_rsci_dinb_d;
  wire [63:0] dout_16_rsci_douta_d;
  wire dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] dout_17_rsci_dinb_d;
  wire [63:0] dout_17_rsci_douta_d;
  wire dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_0_data_rsci_addra_d;
  wire [7:0] tmp_0_data_rsci_addrb_d;
  wire [63:0] tmp_0_data_rsci_dinb_d;
  wire [63:0] tmp_0_data_rsci_douta_d;
  wire tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_1_data_rsci_addra_d;
  wire [7:0] tmp_1_data_rsci_addrb_d;
  wire [63:0] tmp_1_data_rsci_dinb_d;
  wire [63:0] tmp_1_data_rsci_douta_d;
  wire tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_2_data_rsci_addra_d;
  wire [7:0] tmp_2_data_rsci_addrb_d;
  wire [63:0] tmp_2_data_rsci_dinb_d;
  wire [63:0] tmp_2_data_rsci_douta_d;
  wire tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_3_data_rsci_addra_d;
  wire [7:0] tmp_3_data_rsci_addrb_d;
  wire [63:0] tmp_3_data_rsci_dinb_d;
  wire [63:0] tmp_3_data_rsci_douta_d;
  wire tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_4_data_rsci_addra_d;
  wire [7:0] tmp_4_data_rsci_addrb_d;
  wire [63:0] tmp_4_data_rsci_dinb_d;
  wire [63:0] tmp_4_data_rsci_douta_d;
  wire tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_5_data_rsci_addra_d;
  wire [7:0] tmp_5_data_rsci_addrb_d;
  wire [63:0] tmp_5_data_rsci_dinb_d;
  wire [63:0] tmp_5_data_rsci_douta_d;
  wire tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_6_data_rsci_addra_d;
  wire [7:0] tmp_6_data_rsci_addrb_d;
  wire [63:0] tmp_6_data_rsci_dinb_d;
  wire [63:0] tmp_6_data_rsci_douta_d;
  wire tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_7_data_rsci_addra_d;
  wire [7:0] tmp_7_data_rsci_addrb_d;
  wire [63:0] tmp_7_data_rsci_dinb_d;
  wire [63:0] tmp_7_data_rsci_douta_d;
  wire tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_8_data_rsci_addra_d;
  wire [7:0] tmp_8_data_rsci_addrb_d;
  wire [63:0] tmp_8_data_rsci_dinb_d;
  wire [63:0] tmp_8_data_rsci_douta_d;
  wire tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_9_data_rsci_addra_d;
  wire [7:0] tmp_9_data_rsci_addrb_d;
  wire [63:0] tmp_9_data_rsci_dinb_d;
  wire [63:0] tmp_9_data_rsci_douta_d;
  wire tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_10_data_rsci_addra_d;
  wire [7:0] tmp_10_data_rsci_addrb_d;
  wire [63:0] tmp_10_data_rsci_dinb_d;
  wire [63:0] tmp_10_data_rsci_douta_d;
  wire tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_11_data_rsci_addra_d;
  wire [7:0] tmp_11_data_rsci_addrb_d;
  wire [63:0] tmp_11_data_rsci_dinb_d;
  wire [63:0] tmp_11_data_rsci_douta_d;
  wire tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_12_data_rsci_addra_d;
  wire [7:0] tmp_12_data_rsci_addrb_d;
  wire [63:0] tmp_12_data_rsci_dinb_d;
  wire [63:0] tmp_12_data_rsci_douta_d;
  wire tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_13_data_rsci_addra_d;
  wire [7:0] tmp_13_data_rsci_addrb_d;
  wire [63:0] tmp_13_data_rsci_dinb_d;
  wire [63:0] tmp_13_data_rsci_douta_d;
  wire tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_14_data_rsci_addra_d;
  wire [7:0] tmp_14_data_rsci_addrb_d;
  wire [63:0] tmp_14_data_rsci_dinb_d;
  wire [63:0] tmp_14_data_rsci_douta_d;
  wire tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_15_data_rsci_addra_d;
  wire [7:0] tmp_15_data_rsci_addrb_d;
  wire [63:0] tmp_15_data_rsci_dinb_d;
  wire [63:0] tmp_15_data_rsci_douta_d;
  wire tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_16_data_rsci_addra_d;
  wire [7:0] tmp_16_data_rsci_addrb_d;
  wire [63:0] tmp_16_data_rsci_dinb_d;
  wire [63:0] tmp_16_data_rsci_douta_d;
  wire tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] tmp_17_data_rsci_addra_d;
  wire [7:0] tmp_17_data_rsci_addrb_d;
  wire [63:0] tmp_17_data_rsci_dinb_d;
  wire [63:0] tmp_17_data_rsci_douta_d;
  wire tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [63:0] tmp_0_data_rsc_douta;
  wire [63:0] tmp_0_data_rsc_dinb;
  wire [7:0] tmp_0_data_rsc_addrb;
  wire [7:0] tmp_0_data_rsc_addra;
  wire tmp_0_data_rsc_csb_n;
  wire tmp_0_data_rsc_csa_n;
  wire tmp_0_data_rsc_unc_1;
  wire [63:0] tmp_1_data_rsc_douta;
  wire [63:0] tmp_1_data_rsc_dinb;
  wire [7:0] tmp_1_data_rsc_addrb;
  wire [7:0] tmp_1_data_rsc_addra;
  wire tmp_1_data_rsc_csb_n;
  wire tmp_1_data_rsc_csa_n;
  wire tmp_1_data_rsc_unc_1;
  wire [63:0] tmp_2_data_rsc_douta;
  wire [63:0] tmp_2_data_rsc_dinb;
  wire [7:0] tmp_2_data_rsc_addrb;
  wire [7:0] tmp_2_data_rsc_addra;
  wire tmp_2_data_rsc_csb_n;
  wire tmp_2_data_rsc_csa_n;
  wire tmp_2_data_rsc_unc_1;
  wire [63:0] tmp_3_data_rsc_douta;
  wire [63:0] tmp_3_data_rsc_dinb;
  wire [7:0] tmp_3_data_rsc_addrb;
  wire [7:0] tmp_3_data_rsc_addra;
  wire tmp_3_data_rsc_csb_n;
  wire tmp_3_data_rsc_csa_n;
  wire tmp_3_data_rsc_unc_1;
  wire [63:0] tmp_4_data_rsc_douta;
  wire [63:0] tmp_4_data_rsc_dinb;
  wire [7:0] tmp_4_data_rsc_addrb;
  wire [7:0] tmp_4_data_rsc_addra;
  wire tmp_4_data_rsc_csb_n;
  wire tmp_4_data_rsc_csa_n;
  wire tmp_4_data_rsc_unc_1;
  wire [63:0] tmp_5_data_rsc_douta;
  wire [63:0] tmp_5_data_rsc_dinb;
  wire [7:0] tmp_5_data_rsc_addrb;
  wire [7:0] tmp_5_data_rsc_addra;
  wire tmp_5_data_rsc_csb_n;
  wire tmp_5_data_rsc_csa_n;
  wire tmp_5_data_rsc_unc_1;
  wire [63:0] tmp_6_data_rsc_douta;
  wire [63:0] tmp_6_data_rsc_dinb;
  wire [7:0] tmp_6_data_rsc_addrb;
  wire [7:0] tmp_6_data_rsc_addra;
  wire tmp_6_data_rsc_csb_n;
  wire tmp_6_data_rsc_csa_n;
  wire tmp_6_data_rsc_unc_1;
  wire [63:0] tmp_7_data_rsc_douta;
  wire [63:0] tmp_7_data_rsc_dinb;
  wire [7:0] tmp_7_data_rsc_addrb;
  wire [7:0] tmp_7_data_rsc_addra;
  wire tmp_7_data_rsc_csb_n;
  wire tmp_7_data_rsc_csa_n;
  wire tmp_7_data_rsc_unc_1;
  wire [63:0] tmp_8_data_rsc_douta;
  wire [63:0] tmp_8_data_rsc_dinb;
  wire [7:0] tmp_8_data_rsc_addrb;
  wire [7:0] tmp_8_data_rsc_addra;
  wire tmp_8_data_rsc_csb_n;
  wire tmp_8_data_rsc_csa_n;
  wire tmp_8_data_rsc_unc_1;
  wire [63:0] tmp_9_data_rsc_douta;
  wire [63:0] tmp_9_data_rsc_dinb;
  wire [7:0] tmp_9_data_rsc_addrb;
  wire [7:0] tmp_9_data_rsc_addra;
  wire tmp_9_data_rsc_csb_n;
  wire tmp_9_data_rsc_csa_n;
  wire tmp_9_data_rsc_unc_1;
  wire [63:0] tmp_10_data_rsc_douta;
  wire [63:0] tmp_10_data_rsc_dinb;
  wire [7:0] tmp_10_data_rsc_addrb;
  wire [7:0] tmp_10_data_rsc_addra;
  wire tmp_10_data_rsc_csb_n;
  wire tmp_10_data_rsc_csa_n;
  wire tmp_10_data_rsc_unc_1;
  wire [63:0] tmp_11_data_rsc_douta;
  wire [63:0] tmp_11_data_rsc_dinb;
  wire [7:0] tmp_11_data_rsc_addrb;
  wire [7:0] tmp_11_data_rsc_addra;
  wire tmp_11_data_rsc_csb_n;
  wire tmp_11_data_rsc_csa_n;
  wire tmp_11_data_rsc_unc_1;
  wire [63:0] tmp_12_data_rsc_douta;
  wire [63:0] tmp_12_data_rsc_dinb;
  wire [7:0] tmp_12_data_rsc_addrb;
  wire [7:0] tmp_12_data_rsc_addra;
  wire tmp_12_data_rsc_csb_n;
  wire tmp_12_data_rsc_csa_n;
  wire tmp_12_data_rsc_unc_1;
  wire [63:0] tmp_13_data_rsc_douta;
  wire [63:0] tmp_13_data_rsc_dinb;
  wire [7:0] tmp_13_data_rsc_addrb;
  wire [7:0] tmp_13_data_rsc_addra;
  wire tmp_13_data_rsc_csb_n;
  wire tmp_13_data_rsc_csa_n;
  wire tmp_13_data_rsc_unc_1;
  wire [63:0] tmp_14_data_rsc_douta;
  wire [63:0] tmp_14_data_rsc_dinb;
  wire [7:0] tmp_14_data_rsc_addrb;
  wire [7:0] tmp_14_data_rsc_addra;
  wire tmp_14_data_rsc_csb_n;
  wire tmp_14_data_rsc_csa_n;
  wire tmp_14_data_rsc_unc_1;
  wire [63:0] tmp_15_data_rsc_douta;
  wire [63:0] tmp_15_data_rsc_dinb;
  wire [7:0] tmp_15_data_rsc_addrb;
  wire [7:0] tmp_15_data_rsc_addra;
  wire tmp_15_data_rsc_csb_n;
  wire tmp_15_data_rsc_csa_n;
  wire tmp_15_data_rsc_unc_1;
  wire [63:0] tmp_16_data_rsc_douta;
  wire [63:0] tmp_16_data_rsc_dinb;
  wire [7:0] tmp_16_data_rsc_addrb;
  wire [7:0] tmp_16_data_rsc_addra;
  wire tmp_16_data_rsc_csb_n;
  wire tmp_16_data_rsc_csa_n;
  wire tmp_16_data_rsc_unc_1;
  wire [63:0] tmp_17_data_rsc_douta;
  wire [63:0] tmp_17_data_rsc_dinb;
  wire [7:0] tmp_17_data_rsc_addrb;
  wire [7:0] tmp_17_data_rsc_addra;
  wire tmp_17_data_rsc_csb_n;
  wire tmp_17_data_rsc_csa_n;
  wire tmp_17_data_rsc_unc_1;
  wire [6:0] dout_0_rsci_addra_d_iff;
  wire [6:0] dout_1_rsci_addra_d_iff;
  wire [6:0] dout_2_rsci_addra_d_iff;
  wire [6:0] dout_3_rsci_addra_d_iff;
  wire [6:0] dout_4_rsci_addra_d_iff;
  wire [6:0] dout_5_rsci_addra_d_iff;
  wire [6:0] dout_6_rsci_addra_d_iff;
  wire [6:0] dout_7_rsci_addra_d_iff;
  wire [6:0] dout_8_rsci_addra_d_iff;
  wire [6:0] dout_9_rsci_addra_d_iff;
  wire [6:0] dout_10_rsci_addra_d_iff;
  wire [6:0] dout_11_rsci_addra_d_iff;
  wire [6:0] dout_12_rsci_addra_d_iff;
  wire [6:0] dout_13_rsci_addra_d_iff;
  wire [6:0] dout_14_rsci_addra_d_iff;
  wire [6:0] dout_15_rsci_addra_d_iff;
  wire [6:0] dout_16_rsci_addra_d_iff;
  wire [6:0] dout_17_rsci_addra_d_iff;


  // Interconnect Declarations for Component Instantiations 
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_0_data_rsc_comp (
      .addra(tmp_0_data_rsc_addrb),
      .addrb(tmp_0_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_0_data_rsc_csb_n),
      .csb_n(tmp_0_data_rsc_csb_n),
      .dinb(tmp_0_data_rsc_dinb),
      .douta(tmp_0_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_0_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_1_data_rsc_comp (
      .addra(tmp_1_data_rsc_addrb),
      .addrb(tmp_1_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_1_data_rsc_csb_n),
      .csb_n(tmp_1_data_rsc_csb_n),
      .dinb(tmp_1_data_rsc_dinb),
      .douta(tmp_1_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_1_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_2_data_rsc_comp (
      .addra(tmp_2_data_rsc_addrb),
      .addrb(tmp_2_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_2_data_rsc_csb_n),
      .csb_n(tmp_2_data_rsc_csb_n),
      .dinb(tmp_2_data_rsc_dinb),
      .douta(tmp_2_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_2_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_3_data_rsc_comp (
      .addra(tmp_3_data_rsc_addrb),
      .addrb(tmp_3_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_3_data_rsc_csb_n),
      .csb_n(tmp_3_data_rsc_csb_n),
      .dinb(tmp_3_data_rsc_dinb),
      .douta(tmp_3_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_3_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_4_data_rsc_comp (
      .addra(tmp_4_data_rsc_addrb),
      .addrb(tmp_4_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_4_data_rsc_csb_n),
      .csb_n(tmp_4_data_rsc_csb_n),
      .dinb(tmp_4_data_rsc_dinb),
      .douta(tmp_4_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_4_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_5_data_rsc_comp (
      .addra(tmp_5_data_rsc_addrb),
      .addrb(tmp_5_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_5_data_rsc_csb_n),
      .csb_n(tmp_5_data_rsc_csb_n),
      .dinb(tmp_5_data_rsc_dinb),
      .douta(tmp_5_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_5_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_6_data_rsc_comp (
      .addra(tmp_6_data_rsc_addrb),
      .addrb(tmp_6_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_6_data_rsc_csb_n),
      .csb_n(tmp_6_data_rsc_csb_n),
      .dinb(tmp_6_data_rsc_dinb),
      .douta(tmp_6_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_6_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_7_data_rsc_comp (
      .addra(tmp_7_data_rsc_addrb),
      .addrb(tmp_7_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_7_data_rsc_csb_n),
      .csb_n(tmp_7_data_rsc_csb_n),
      .dinb(tmp_7_data_rsc_dinb),
      .douta(tmp_7_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_7_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_8_data_rsc_comp (
      .addra(tmp_8_data_rsc_addrb),
      .addrb(tmp_8_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_8_data_rsc_csb_n),
      .csb_n(tmp_8_data_rsc_csb_n),
      .dinb(tmp_8_data_rsc_dinb),
      .douta(tmp_8_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_8_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_9_data_rsc_comp (
      .addra(tmp_9_data_rsc_addrb),
      .addrb(tmp_9_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_9_data_rsc_csb_n),
      .csb_n(tmp_9_data_rsc_csb_n),
      .dinb(tmp_9_data_rsc_dinb),
      .douta(tmp_9_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_9_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_10_data_rsc_comp (
      .addra(tmp_10_data_rsc_addrb),
      .addrb(tmp_10_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_10_data_rsc_csb_n),
      .csb_n(tmp_10_data_rsc_csb_n),
      .dinb(tmp_10_data_rsc_dinb),
      .douta(tmp_10_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_10_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_11_data_rsc_comp (
      .addra(tmp_11_data_rsc_addrb),
      .addrb(tmp_11_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_11_data_rsc_csb_n),
      .csb_n(tmp_11_data_rsc_csb_n),
      .dinb(tmp_11_data_rsc_dinb),
      .douta(tmp_11_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_11_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_12_data_rsc_comp (
      .addra(tmp_12_data_rsc_addrb),
      .addrb(tmp_12_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_12_data_rsc_csb_n),
      .csb_n(tmp_12_data_rsc_csb_n),
      .dinb(tmp_12_data_rsc_dinb),
      .douta(tmp_12_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_12_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_13_data_rsc_comp (
      .addra(tmp_13_data_rsc_addrb),
      .addrb(tmp_13_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_13_data_rsc_csb_n),
      .csb_n(tmp_13_data_rsc_csb_n),
      .dinb(tmp_13_data_rsc_dinb),
      .douta(tmp_13_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_13_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_14_data_rsc_comp (
      .addra(tmp_14_data_rsc_addrb),
      .addrb(tmp_14_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_14_data_rsc_csb_n),
      .csb_n(tmp_14_data_rsc_csb_n),
      .dinb(tmp_14_data_rsc_dinb),
      .douta(tmp_14_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_14_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_15_data_rsc_comp (
      .addra(tmp_15_data_rsc_addrb),
      .addrb(tmp_15_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_15_data_rsc_csb_n),
      .csb_n(tmp_15_data_rsc_csb_n),
      .dinb(tmp_15_data_rsc_dinb),
      .douta(tmp_15_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_15_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_16_data_rsc_comp (
      .addra(tmp_16_data_rsc_addrb),
      .addrb(tmp_16_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_16_data_rsc_csb_n),
      .csb_n(tmp_16_data_rsc_csb_n),
      .dinb(tmp_16_data_rsc_dinb),
      .douta(tmp_16_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_16_data_rsc_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) tmp_17_data_rsc_comp (
      .addra(tmp_17_data_rsc_addrb),
      .addrb(tmp_17_data_rsc_addrb),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(tmp_17_data_rsc_csb_n),
      .csb_n(tmp_17_data_rsc_csb_n),
      .dinb(tmp_17_data_rsc_dinb),
      .douta(tmp_17_data_rsc_douta),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(tmp_17_data_rsc_unc_1)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_2_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_0_rsci (
      .douta(dout_0_rsc_douta),
      .dinb(dout_0_rsc_dinb),
      .addrb(dout_0_rsc_addrb),
      .addra(dout_0_rsc_addra),
      .csb_n(dout_0_rsc_csb_n),
      .csa_n(dout_0_rsc_csa_n),
      .addra_d(dout_0_rsci_addra_d_iff),
      .addrb_d(dout_0_rsci_addra_d_iff),
      .dinb_d(dout_0_rsci_dinb_d),
      .douta_d(dout_0_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_3_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_1_rsci (
      .douta(dout_1_rsc_douta),
      .dinb(dout_1_rsc_dinb),
      .addrb(dout_1_rsc_addrb),
      .addra(dout_1_rsc_addra),
      .csb_n(dout_1_rsc_csb_n),
      .csa_n(dout_1_rsc_csa_n),
      .addra_d(dout_1_rsci_addra_d_iff),
      .addrb_d(dout_1_rsci_addra_d_iff),
      .dinb_d(dout_1_rsci_dinb_d),
      .douta_d(dout_1_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_4_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_2_rsci (
      .douta(dout_2_rsc_douta),
      .dinb(dout_2_rsc_dinb),
      .addrb(dout_2_rsc_addrb),
      .addra(dout_2_rsc_addra),
      .csb_n(dout_2_rsc_csb_n),
      .csa_n(dout_2_rsc_csa_n),
      .addra_d(dout_2_rsci_addra_d_iff),
      .addrb_d(dout_2_rsci_addra_d_iff),
      .dinb_d(dout_2_rsci_dinb_d),
      .douta_d(dout_2_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_5_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_3_rsci (
      .douta(dout_3_rsc_douta),
      .dinb(dout_3_rsc_dinb),
      .addrb(dout_3_rsc_addrb),
      .addra(dout_3_rsc_addra),
      .csb_n(dout_3_rsc_csb_n),
      .csa_n(dout_3_rsc_csa_n),
      .addra_d(dout_3_rsci_addra_d_iff),
      .addrb_d(dout_3_rsci_addra_d_iff),
      .dinb_d(dout_3_rsci_dinb_d),
      .douta_d(dout_3_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_6_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_4_rsci (
      .douta(dout_4_rsc_douta),
      .dinb(dout_4_rsc_dinb),
      .addrb(dout_4_rsc_addrb),
      .addra(dout_4_rsc_addra),
      .csb_n(dout_4_rsc_csb_n),
      .csa_n(dout_4_rsc_csa_n),
      .addra_d(dout_4_rsci_addra_d_iff),
      .addrb_d(dout_4_rsci_addra_d_iff),
      .dinb_d(dout_4_rsci_dinb_d),
      .douta_d(dout_4_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_7_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_5_rsci (
      .douta(dout_5_rsc_douta),
      .dinb(dout_5_rsc_dinb),
      .addrb(dout_5_rsc_addrb),
      .addra(dout_5_rsc_addra),
      .csb_n(dout_5_rsc_csb_n),
      .csa_n(dout_5_rsc_csa_n),
      .addra_d(dout_5_rsci_addra_d_iff),
      .addrb_d(dout_5_rsci_addra_d_iff),
      .dinb_d(dout_5_rsci_dinb_d),
      .douta_d(dout_5_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_8_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_6_rsci (
      .douta(dout_6_rsc_douta),
      .dinb(dout_6_rsc_dinb),
      .addrb(dout_6_rsc_addrb),
      .addra(dout_6_rsc_addra),
      .csb_n(dout_6_rsc_csb_n),
      .csa_n(dout_6_rsc_csa_n),
      .addra_d(dout_6_rsci_addra_d_iff),
      .addrb_d(dout_6_rsci_addra_d_iff),
      .dinb_d(dout_6_rsci_dinb_d),
      .douta_d(dout_6_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_9_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_7_rsci (
      .douta(dout_7_rsc_douta),
      .dinb(dout_7_rsc_dinb),
      .addrb(dout_7_rsc_addrb),
      .addra(dout_7_rsc_addra),
      .csb_n(dout_7_rsc_csb_n),
      .csa_n(dout_7_rsc_csa_n),
      .addra_d(dout_7_rsci_addra_d_iff),
      .addrb_d(dout_7_rsci_addra_d_iff),
      .dinb_d(dout_7_rsci_dinb_d),
      .douta_d(dout_7_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_10_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_8_rsci (
      .douta(dout_8_rsc_douta),
      .dinb(dout_8_rsc_dinb),
      .addrb(dout_8_rsc_addrb),
      .addra(dout_8_rsc_addra),
      .csb_n(dout_8_rsc_csb_n),
      .csa_n(dout_8_rsc_csa_n),
      .addra_d(dout_8_rsci_addra_d_iff),
      .addrb_d(dout_8_rsci_addra_d_iff),
      .dinb_d(dout_8_rsci_dinb_d),
      .douta_d(dout_8_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_11_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_9_rsci (
      .douta(dout_9_rsc_douta),
      .dinb(dout_9_rsc_dinb),
      .addrb(dout_9_rsc_addrb),
      .addra(dout_9_rsc_addra),
      .csb_n(dout_9_rsc_csb_n),
      .csa_n(dout_9_rsc_csa_n),
      .addra_d(dout_9_rsci_addra_d_iff),
      .addrb_d(dout_9_rsci_addra_d_iff),
      .dinb_d(dout_9_rsci_dinb_d),
      .douta_d(dout_9_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_12_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_10_rsci (
      .douta(dout_10_rsc_douta),
      .dinb(dout_10_rsc_dinb),
      .addrb(dout_10_rsc_addrb),
      .addra(dout_10_rsc_addra),
      .csb_n(dout_10_rsc_csb_n),
      .csa_n(dout_10_rsc_csa_n),
      .addra_d(dout_10_rsci_addra_d_iff),
      .addrb_d(dout_10_rsci_addra_d_iff),
      .dinb_d(dout_10_rsci_dinb_d),
      .douta_d(dout_10_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_13_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_11_rsci (
      .douta(dout_11_rsc_douta),
      .dinb(dout_11_rsc_dinb),
      .addrb(dout_11_rsc_addrb),
      .addra(dout_11_rsc_addra),
      .csb_n(dout_11_rsc_csb_n),
      .csa_n(dout_11_rsc_csa_n),
      .addra_d(dout_11_rsci_addra_d_iff),
      .addrb_d(dout_11_rsci_addra_d_iff),
      .dinb_d(dout_11_rsci_dinb_d),
      .douta_d(dout_11_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_14_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_12_rsci (
      .douta(dout_12_rsc_douta),
      .dinb(dout_12_rsc_dinb),
      .addrb(dout_12_rsc_addrb),
      .addra(dout_12_rsc_addra),
      .csb_n(dout_12_rsc_csb_n),
      .csa_n(dout_12_rsc_csa_n),
      .addra_d(dout_12_rsci_addra_d_iff),
      .addrb_d(dout_12_rsci_addra_d_iff),
      .dinb_d(dout_12_rsci_dinb_d),
      .douta_d(dout_12_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_15_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_13_rsci (
      .douta(dout_13_rsc_douta),
      .dinb(dout_13_rsc_dinb),
      .addrb(dout_13_rsc_addrb),
      .addra(dout_13_rsc_addra),
      .csb_n(dout_13_rsc_csb_n),
      .csa_n(dout_13_rsc_csa_n),
      .addra_d(dout_13_rsci_addra_d_iff),
      .addrb_d(dout_13_rsci_addra_d_iff),
      .dinb_d(dout_13_rsci_dinb_d),
      .douta_d(dout_13_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_16_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_14_rsci (
      .douta(dout_14_rsc_douta),
      .dinb(dout_14_rsc_dinb),
      .addrb(dout_14_rsc_addrb),
      .addra(dout_14_rsc_addra),
      .csb_n(dout_14_rsc_csb_n),
      .csa_n(dout_14_rsc_csa_n),
      .addra_d(dout_14_rsci_addra_d_iff),
      .addrb_d(dout_14_rsci_addra_d_iff),
      .dinb_d(dout_14_rsci_dinb_d),
      .douta_d(dout_14_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_17_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_15_rsci (
      .douta(dout_15_rsc_douta),
      .dinb(dout_15_rsc_dinb),
      .addrb(dout_15_rsc_addrb),
      .addra(dout_15_rsc_addra),
      .csb_n(dout_15_rsc_csb_n),
      .csa_n(dout_15_rsc_csa_n),
      .addra_d(dout_15_rsci_addra_d_iff),
      .addrb_d(dout_15_rsci_addra_d_iff),
      .dinb_d(dout_15_rsci_dinb_d),
      .douta_d(dout_15_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_18_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_16_rsci (
      .douta(dout_16_rsc_douta),
      .dinb(dout_16_rsc_dinb),
      .addrb(dout_16_rsc_addrb),
      .addra(dout_16_rsc_addra),
      .csb_n(dout_16_rsc_csb_n),
      .csa_n(dout_16_rsc_csa_n),
      .addra_d(dout_16_rsci_addra_d_iff),
      .addrb_d(dout_16_rsci_addra_d_iff),
      .dinb_d(dout_16_rsci_dinb_d),
      .douta_d(dout_16_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_19_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      dout_17_rsci (
      .douta(dout_17_rsc_douta),
      .dinb(dout_17_rsc_dinb),
      .addrb(dout_17_rsc_addrb),
      .addra(dout_17_rsc_addra),
      .csb_n(dout_17_rsc_csb_n),
      .csa_n(dout_17_rsc_csa_n),
      .addra_d(dout_17_rsci_addra_d_iff),
      .addrb_d(dout_17_rsci_addra_d_iff),
      .dinb_d(dout_17_rsci_dinb_d),
      .douta_d(dout_17_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_20_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_0_data_rsci (
      .douta(tmp_0_data_rsc_douta),
      .dinb(tmp_0_data_rsc_dinb),
      .addrb(tmp_0_data_rsc_addrb),
      .addra(tmp_0_data_rsc_addra),
      .csb_n(tmp_0_data_rsc_csb_n),
      .csa_n(tmp_0_data_rsc_csa_n),
      .addra_d(tmp_0_data_rsci_addra_d),
      .addrb_d(tmp_0_data_rsci_addrb_d),
      .dinb_d(tmp_0_data_rsci_dinb_d),
      .douta_d(tmp_0_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_21_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_1_data_rsci (
      .douta(tmp_1_data_rsc_douta),
      .dinb(tmp_1_data_rsc_dinb),
      .addrb(tmp_1_data_rsc_addrb),
      .addra(tmp_1_data_rsc_addra),
      .csb_n(tmp_1_data_rsc_csb_n),
      .csa_n(tmp_1_data_rsc_csa_n),
      .addra_d(tmp_1_data_rsci_addra_d),
      .addrb_d(tmp_1_data_rsci_addrb_d),
      .dinb_d(tmp_1_data_rsci_dinb_d),
      .douta_d(tmp_1_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_22_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_2_data_rsci (
      .douta(tmp_2_data_rsc_douta),
      .dinb(tmp_2_data_rsc_dinb),
      .addrb(tmp_2_data_rsc_addrb),
      .addra(tmp_2_data_rsc_addra),
      .csb_n(tmp_2_data_rsc_csb_n),
      .csa_n(tmp_2_data_rsc_csa_n),
      .addra_d(tmp_2_data_rsci_addra_d),
      .addrb_d(tmp_2_data_rsci_addrb_d),
      .dinb_d(tmp_2_data_rsci_dinb_d),
      .douta_d(tmp_2_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_23_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_3_data_rsci (
      .douta(tmp_3_data_rsc_douta),
      .dinb(tmp_3_data_rsc_dinb),
      .addrb(tmp_3_data_rsc_addrb),
      .addra(tmp_3_data_rsc_addra),
      .csb_n(tmp_3_data_rsc_csb_n),
      .csa_n(tmp_3_data_rsc_csa_n),
      .addra_d(tmp_3_data_rsci_addra_d),
      .addrb_d(tmp_3_data_rsci_addrb_d),
      .dinb_d(tmp_3_data_rsci_dinb_d),
      .douta_d(tmp_3_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_24_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_4_data_rsci (
      .douta(tmp_4_data_rsc_douta),
      .dinb(tmp_4_data_rsc_dinb),
      .addrb(tmp_4_data_rsc_addrb),
      .addra(tmp_4_data_rsc_addra),
      .csb_n(tmp_4_data_rsc_csb_n),
      .csa_n(tmp_4_data_rsc_csa_n),
      .addra_d(tmp_4_data_rsci_addra_d),
      .addrb_d(tmp_4_data_rsci_addrb_d),
      .dinb_d(tmp_4_data_rsci_dinb_d),
      .douta_d(tmp_4_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_25_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_5_data_rsci (
      .douta(tmp_5_data_rsc_douta),
      .dinb(tmp_5_data_rsc_dinb),
      .addrb(tmp_5_data_rsc_addrb),
      .addra(tmp_5_data_rsc_addra),
      .csb_n(tmp_5_data_rsc_csb_n),
      .csa_n(tmp_5_data_rsc_csa_n),
      .addra_d(tmp_5_data_rsci_addra_d),
      .addrb_d(tmp_5_data_rsci_addrb_d),
      .dinb_d(tmp_5_data_rsci_dinb_d),
      .douta_d(tmp_5_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_26_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_6_data_rsci (
      .douta(tmp_6_data_rsc_douta),
      .dinb(tmp_6_data_rsc_dinb),
      .addrb(tmp_6_data_rsc_addrb),
      .addra(tmp_6_data_rsc_addra),
      .csb_n(tmp_6_data_rsc_csb_n),
      .csa_n(tmp_6_data_rsc_csa_n),
      .addra_d(tmp_6_data_rsci_addra_d),
      .addrb_d(tmp_6_data_rsci_addrb_d),
      .dinb_d(tmp_6_data_rsci_dinb_d),
      .douta_d(tmp_6_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_27_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_7_data_rsci (
      .douta(tmp_7_data_rsc_douta),
      .dinb(tmp_7_data_rsc_dinb),
      .addrb(tmp_7_data_rsc_addrb),
      .addra(tmp_7_data_rsc_addra),
      .csb_n(tmp_7_data_rsc_csb_n),
      .csa_n(tmp_7_data_rsc_csa_n),
      .addra_d(tmp_7_data_rsci_addra_d),
      .addrb_d(tmp_7_data_rsci_addrb_d),
      .dinb_d(tmp_7_data_rsci_dinb_d),
      .douta_d(tmp_7_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_28_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_8_data_rsci (
      .douta(tmp_8_data_rsc_douta),
      .dinb(tmp_8_data_rsc_dinb),
      .addrb(tmp_8_data_rsc_addrb),
      .addra(tmp_8_data_rsc_addra),
      .csb_n(tmp_8_data_rsc_csb_n),
      .csa_n(tmp_8_data_rsc_csa_n),
      .addra_d(tmp_8_data_rsci_addra_d),
      .addrb_d(tmp_8_data_rsci_addrb_d),
      .dinb_d(tmp_8_data_rsci_dinb_d),
      .douta_d(tmp_8_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_29_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_9_data_rsci (
      .douta(tmp_9_data_rsc_douta),
      .dinb(tmp_9_data_rsc_dinb),
      .addrb(tmp_9_data_rsc_addrb),
      .addra(tmp_9_data_rsc_addra),
      .csb_n(tmp_9_data_rsc_csb_n),
      .csa_n(tmp_9_data_rsc_csa_n),
      .addra_d(tmp_9_data_rsci_addra_d),
      .addrb_d(tmp_9_data_rsci_addrb_d),
      .dinb_d(tmp_9_data_rsci_dinb_d),
      .douta_d(tmp_9_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_30_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_10_data_rsci (
      .douta(tmp_10_data_rsc_douta),
      .dinb(tmp_10_data_rsc_dinb),
      .addrb(tmp_10_data_rsc_addrb),
      .addra(tmp_10_data_rsc_addra),
      .csb_n(tmp_10_data_rsc_csb_n),
      .csa_n(tmp_10_data_rsc_csa_n),
      .addra_d(tmp_10_data_rsci_addra_d),
      .addrb_d(tmp_10_data_rsci_addrb_d),
      .dinb_d(tmp_10_data_rsci_dinb_d),
      .douta_d(tmp_10_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_31_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_11_data_rsci (
      .douta(tmp_11_data_rsc_douta),
      .dinb(tmp_11_data_rsc_dinb),
      .addrb(tmp_11_data_rsc_addrb),
      .addra(tmp_11_data_rsc_addra),
      .csb_n(tmp_11_data_rsc_csb_n),
      .csa_n(tmp_11_data_rsc_csa_n),
      .addra_d(tmp_11_data_rsci_addra_d),
      .addrb_d(tmp_11_data_rsci_addrb_d),
      .dinb_d(tmp_11_data_rsci_dinb_d),
      .douta_d(tmp_11_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_32_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_12_data_rsci (
      .douta(tmp_12_data_rsc_douta),
      .dinb(tmp_12_data_rsc_dinb),
      .addrb(tmp_12_data_rsc_addrb),
      .addra(tmp_12_data_rsc_addra),
      .csb_n(tmp_12_data_rsc_csb_n),
      .csa_n(tmp_12_data_rsc_csa_n),
      .addra_d(tmp_12_data_rsci_addra_d),
      .addrb_d(tmp_12_data_rsci_addrb_d),
      .dinb_d(tmp_12_data_rsci_dinb_d),
      .douta_d(tmp_12_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_33_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_13_data_rsci (
      .douta(tmp_13_data_rsc_douta),
      .dinb(tmp_13_data_rsc_dinb),
      .addrb(tmp_13_data_rsc_addrb),
      .addra(tmp_13_data_rsc_addra),
      .csb_n(tmp_13_data_rsc_csb_n),
      .csa_n(tmp_13_data_rsc_csa_n),
      .addra_d(tmp_13_data_rsci_addra_d),
      .addrb_d(tmp_13_data_rsci_addrb_d),
      .dinb_d(tmp_13_data_rsci_dinb_d),
      .douta_d(tmp_13_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_34_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_14_data_rsci (
      .douta(tmp_14_data_rsc_douta),
      .dinb(tmp_14_data_rsc_dinb),
      .addrb(tmp_14_data_rsc_addrb),
      .addra(tmp_14_data_rsc_addra),
      .csb_n(tmp_14_data_rsc_csb_n),
      .csa_n(tmp_14_data_rsc_csa_n),
      .addra_d(tmp_14_data_rsci_addra_d),
      .addrb_d(tmp_14_data_rsci_addrb_d),
      .dinb_d(tmp_14_data_rsci_dinb_d),
      .douta_d(tmp_14_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_35_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_15_data_rsci (
      .douta(tmp_15_data_rsc_douta),
      .dinb(tmp_15_data_rsc_dinb),
      .addrb(tmp_15_data_rsc_addrb),
      .addra(tmp_15_data_rsc_addra),
      .csb_n(tmp_15_data_rsc_csb_n),
      .csa_n(tmp_15_data_rsc_csa_n),
      .addra_d(tmp_15_data_rsci_addra_d),
      .addrb_d(tmp_15_data_rsci_addrb_d),
      .dinb_d(tmp_15_data_rsci_dinb_d),
      .douta_d(tmp_15_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_36_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_16_data_rsci (
      .douta(tmp_16_data_rsc_douta),
      .dinb(tmp_16_data_rsc_dinb),
      .addrb(tmp_16_data_rsc_addrb),
      .addra(tmp_16_data_rsc_addra),
      .csb_n(tmp_16_data_rsc_csb_n),
      .csa_n(tmp_16_data_rsc_csa_n),
      .addra_d(tmp_16_data_rsci_addra_d),
      .addrb_d(tmp_16_data_rsci_addrb_d),
      .dinb_d(tmp_16_data_rsci_dinb_d),
      .douta_d(tmp_16_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_37_n1073741823_n1073741823_66_16_256_0_0_0_0_0_0_0_gen
      tmp_17_data_rsci (
      .douta(tmp_17_data_rsc_douta),
      .dinb(tmp_17_data_rsc_dinb),
      .addrb(tmp_17_data_rsc_addrb),
      .addra(tmp_17_data_rsc_addra),
      .csb_n(tmp_17_data_rsc_csb_n),
      .csa_n(tmp_17_data_rsc_csa_n),
      .addra_d(tmp_17_data_rsci_addra_d),
      .addrb_d(tmp_17_data_rsci_addrb_d),
      .dinb_d(tmp_17_data_rsci_dinb_d),
      .douta_d(tmp_17_data_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_core_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(din_rsc_z),
      .din_rsc_vz(din_rsc_vz),
      .din_rsc_lz(din_rsc_lz),
      .dout_0_rsc_req_vz(dout_0_rsc_req_vz),
      .dout_0_rsc_rls_lz(dout_0_rsc_rls_lz),
      .dout_1_rsc_req_vz(dout_1_rsc_req_vz),
      .dout_1_rsc_rls_lz(dout_1_rsc_rls_lz),
      .dout_2_rsc_req_vz(dout_2_rsc_req_vz),
      .dout_2_rsc_rls_lz(dout_2_rsc_rls_lz),
      .dout_3_rsc_req_vz(dout_3_rsc_req_vz),
      .dout_3_rsc_rls_lz(dout_3_rsc_rls_lz),
      .dout_4_rsc_req_vz(dout_4_rsc_req_vz),
      .dout_4_rsc_rls_lz(dout_4_rsc_rls_lz),
      .dout_5_rsc_req_vz(dout_5_rsc_req_vz),
      .dout_5_rsc_rls_lz(dout_5_rsc_rls_lz),
      .dout_6_rsc_req_vz(dout_6_rsc_req_vz),
      .dout_6_rsc_rls_lz(dout_6_rsc_rls_lz),
      .dout_7_rsc_req_vz(dout_7_rsc_req_vz),
      .dout_7_rsc_rls_lz(dout_7_rsc_rls_lz),
      .dout_8_rsc_req_vz(dout_8_rsc_req_vz),
      .dout_8_rsc_rls_lz(dout_8_rsc_rls_lz),
      .dout_9_rsc_req_vz(dout_9_rsc_req_vz),
      .dout_9_rsc_rls_lz(dout_9_rsc_rls_lz),
      .dout_10_rsc_req_vz(dout_10_rsc_req_vz),
      .dout_10_rsc_rls_lz(dout_10_rsc_rls_lz),
      .dout_11_rsc_req_vz(dout_11_rsc_req_vz),
      .dout_11_rsc_rls_lz(dout_11_rsc_rls_lz),
      .dout_12_rsc_req_vz(dout_12_rsc_req_vz),
      .dout_12_rsc_rls_lz(dout_12_rsc_rls_lz),
      .dout_13_rsc_req_vz(dout_13_rsc_req_vz),
      .dout_13_rsc_rls_lz(dout_13_rsc_rls_lz),
      .dout_14_rsc_req_vz(dout_14_rsc_req_vz),
      .dout_14_rsc_rls_lz(dout_14_rsc_rls_lz),
      .dout_15_rsc_req_vz(dout_15_rsc_req_vz),
      .dout_15_rsc_rls_lz(dout_15_rsc_rls_lz),
      .dout_16_rsc_req_vz(dout_16_rsc_req_vz),
      .dout_16_rsc_rls_lz(dout_16_rsc_rls_lz),
      .dout_17_rsc_req_vz(dout_17_rsc_req_vz),
      .dout_17_rsc_rls_lz(dout_17_rsc_rls_lz),
      .dout_0_rsci_dinb_d(dout_0_rsci_dinb_d),
      .dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_1_rsci_dinb_d(dout_1_rsci_dinb_d),
      .dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_2_rsci_dinb_d(dout_2_rsci_dinb_d),
      .dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_3_rsci_dinb_d(dout_3_rsci_dinb_d),
      .dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_4_rsci_dinb_d(dout_4_rsci_dinb_d),
      .dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_5_rsci_dinb_d(dout_5_rsci_dinb_d),
      .dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_6_rsci_dinb_d(dout_6_rsci_dinb_d),
      .dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_7_rsci_dinb_d(dout_7_rsci_dinb_d),
      .dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_8_rsci_dinb_d(dout_8_rsci_dinb_d),
      .dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_9_rsci_dinb_d(dout_9_rsci_dinb_d),
      .dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_10_rsci_dinb_d(dout_10_rsci_dinb_d),
      .dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_11_rsci_dinb_d(dout_11_rsci_dinb_d),
      .dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_12_rsci_dinb_d(dout_12_rsci_dinb_d),
      .dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_13_rsci_dinb_d(dout_13_rsci_dinb_d),
      .dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_14_rsci_dinb_d(dout_14_rsci_dinb_d),
      .dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_15_rsci_dinb_d(dout_15_rsci_dinb_d),
      .dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_16_rsci_dinb_d(dout_16_rsci_dinb_d),
      .dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_16_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_17_rsci_dinb_d(dout_17_rsci_dinb_d),
      .dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_17_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_0_data_rsci_addra_d(tmp_0_data_rsci_addra_d),
      .tmp_0_data_rsci_addrb_d(tmp_0_data_rsci_addrb_d),
      .tmp_0_data_rsci_dinb_d(tmp_0_data_rsci_dinb_d),
      .tmp_0_data_rsci_douta_d(tmp_0_data_rsci_douta_d),
      .tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_0_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_0_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_1_data_rsci_addra_d(tmp_1_data_rsci_addra_d),
      .tmp_1_data_rsci_addrb_d(tmp_1_data_rsci_addrb_d),
      .tmp_1_data_rsci_dinb_d(tmp_1_data_rsci_dinb_d),
      .tmp_1_data_rsci_douta_d(tmp_1_data_rsci_douta_d),
      .tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_1_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_1_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_2_data_rsci_addra_d(tmp_2_data_rsci_addra_d),
      .tmp_2_data_rsci_addrb_d(tmp_2_data_rsci_addrb_d),
      .tmp_2_data_rsci_dinb_d(tmp_2_data_rsci_dinb_d),
      .tmp_2_data_rsci_douta_d(tmp_2_data_rsci_douta_d),
      .tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_2_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_2_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_3_data_rsci_addra_d(tmp_3_data_rsci_addra_d),
      .tmp_3_data_rsci_addrb_d(tmp_3_data_rsci_addrb_d),
      .tmp_3_data_rsci_dinb_d(tmp_3_data_rsci_dinb_d),
      .tmp_3_data_rsci_douta_d(tmp_3_data_rsci_douta_d),
      .tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_3_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_3_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_4_data_rsci_addra_d(tmp_4_data_rsci_addra_d),
      .tmp_4_data_rsci_addrb_d(tmp_4_data_rsci_addrb_d),
      .tmp_4_data_rsci_dinb_d(tmp_4_data_rsci_dinb_d),
      .tmp_4_data_rsci_douta_d(tmp_4_data_rsci_douta_d),
      .tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_4_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_4_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_5_data_rsci_addra_d(tmp_5_data_rsci_addra_d),
      .tmp_5_data_rsci_addrb_d(tmp_5_data_rsci_addrb_d),
      .tmp_5_data_rsci_dinb_d(tmp_5_data_rsci_dinb_d),
      .tmp_5_data_rsci_douta_d(tmp_5_data_rsci_douta_d),
      .tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_5_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_5_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_6_data_rsci_addra_d(tmp_6_data_rsci_addra_d),
      .tmp_6_data_rsci_addrb_d(tmp_6_data_rsci_addrb_d),
      .tmp_6_data_rsci_dinb_d(tmp_6_data_rsci_dinb_d),
      .tmp_6_data_rsci_douta_d(tmp_6_data_rsci_douta_d),
      .tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_6_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_6_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_7_data_rsci_addra_d(tmp_7_data_rsci_addra_d),
      .tmp_7_data_rsci_addrb_d(tmp_7_data_rsci_addrb_d),
      .tmp_7_data_rsci_dinb_d(tmp_7_data_rsci_dinb_d),
      .tmp_7_data_rsci_douta_d(tmp_7_data_rsci_douta_d),
      .tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_7_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_7_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_8_data_rsci_addra_d(tmp_8_data_rsci_addra_d),
      .tmp_8_data_rsci_addrb_d(tmp_8_data_rsci_addrb_d),
      .tmp_8_data_rsci_dinb_d(tmp_8_data_rsci_dinb_d),
      .tmp_8_data_rsci_douta_d(tmp_8_data_rsci_douta_d),
      .tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_8_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_8_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_9_data_rsci_addra_d(tmp_9_data_rsci_addra_d),
      .tmp_9_data_rsci_addrb_d(tmp_9_data_rsci_addrb_d),
      .tmp_9_data_rsci_dinb_d(tmp_9_data_rsci_dinb_d),
      .tmp_9_data_rsci_douta_d(tmp_9_data_rsci_douta_d),
      .tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_9_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_9_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_10_data_rsci_addra_d(tmp_10_data_rsci_addra_d),
      .tmp_10_data_rsci_addrb_d(tmp_10_data_rsci_addrb_d),
      .tmp_10_data_rsci_dinb_d(tmp_10_data_rsci_dinb_d),
      .tmp_10_data_rsci_douta_d(tmp_10_data_rsci_douta_d),
      .tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_10_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_10_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_11_data_rsci_addra_d(tmp_11_data_rsci_addra_d),
      .tmp_11_data_rsci_addrb_d(tmp_11_data_rsci_addrb_d),
      .tmp_11_data_rsci_dinb_d(tmp_11_data_rsci_dinb_d),
      .tmp_11_data_rsci_douta_d(tmp_11_data_rsci_douta_d),
      .tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_11_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_11_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_12_data_rsci_addra_d(tmp_12_data_rsci_addra_d),
      .tmp_12_data_rsci_addrb_d(tmp_12_data_rsci_addrb_d),
      .tmp_12_data_rsci_dinb_d(tmp_12_data_rsci_dinb_d),
      .tmp_12_data_rsci_douta_d(tmp_12_data_rsci_douta_d),
      .tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_12_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_12_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_13_data_rsci_addra_d(tmp_13_data_rsci_addra_d),
      .tmp_13_data_rsci_addrb_d(tmp_13_data_rsci_addrb_d),
      .tmp_13_data_rsci_dinb_d(tmp_13_data_rsci_dinb_d),
      .tmp_13_data_rsci_douta_d(tmp_13_data_rsci_douta_d),
      .tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_13_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_13_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_14_data_rsci_addra_d(tmp_14_data_rsci_addra_d),
      .tmp_14_data_rsci_addrb_d(tmp_14_data_rsci_addrb_d),
      .tmp_14_data_rsci_dinb_d(tmp_14_data_rsci_dinb_d),
      .tmp_14_data_rsci_douta_d(tmp_14_data_rsci_douta_d),
      .tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_14_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_14_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_15_data_rsci_addra_d(tmp_15_data_rsci_addra_d),
      .tmp_15_data_rsci_addrb_d(tmp_15_data_rsci_addrb_d),
      .tmp_15_data_rsci_dinb_d(tmp_15_data_rsci_dinb_d),
      .tmp_15_data_rsci_douta_d(tmp_15_data_rsci_douta_d),
      .tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_15_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_15_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_16_data_rsci_addra_d(tmp_16_data_rsci_addra_d),
      .tmp_16_data_rsci_addrb_d(tmp_16_data_rsci_addrb_d),
      .tmp_16_data_rsci_dinb_d(tmp_16_data_rsci_dinb_d),
      .tmp_16_data_rsci_douta_d(tmp_16_data_rsci_douta_d),
      .tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_16_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_16_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .tmp_17_data_rsci_addra_d(tmp_17_data_rsci_addra_d),
      .tmp_17_data_rsci_addrb_d(tmp_17_data_rsci_addrb_d),
      .tmp_17_data_rsci_dinb_d(tmp_17_data_rsci_dinb_d),
      .tmp_17_data_rsci_douta_d(tmp_17_data_rsci_douta_d),
      .tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(tmp_17_data_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(tmp_17_data_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_0_rsci_addra_d_pff(dout_0_rsci_addra_d_iff),
      .dout_1_rsci_addra_d_pff(dout_1_rsci_addra_d_iff),
      .dout_2_rsci_addra_d_pff(dout_2_rsci_addra_d_iff),
      .dout_3_rsci_addra_d_pff(dout_3_rsci_addra_d_iff),
      .dout_4_rsci_addra_d_pff(dout_4_rsci_addra_d_iff),
      .dout_5_rsci_addra_d_pff(dout_5_rsci_addra_d_iff),
      .dout_6_rsci_addra_d_pff(dout_6_rsci_addra_d_iff),
      .dout_7_rsci_addra_d_pff(dout_7_rsci_addra_d_iff),
      .dout_8_rsci_addra_d_pff(dout_8_rsci_addra_d_iff),
      .dout_9_rsci_addra_d_pff(dout_9_rsci_addra_d_iff),
      .dout_10_rsci_addra_d_pff(dout_10_rsci_addra_d_iff),
      .dout_11_rsci_addra_d_pff(dout_11_rsci_addra_d_iff),
      .dout_12_rsci_addra_d_pff(dout_12_rsci_addra_d_iff),
      .dout_13_rsci_addra_d_pff(dout_13_rsci_addra_d_iff),
      .dout_14_rsci_addra_d_pff(dout_14_rsci_addra_d_iff),
      .dout_15_rsci_addra_d_pff(dout_15_rsci_addra_d_iff),
      .dout_16_rsci_addra_d_pff(dout_16_rsci_addra_d_iff),
      .dout_17_rsci_addra_d_pff(dout_17_rsci_addra_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_1
// ------------------------------------------------------------------


module READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_1 (
  clk, rst, din_0_rsc_csa_n, din_0_rsc_csb_n, din_0_rsc_addra, din_0_rsc_addrb, din_0_rsc_dinb,
      din_0_rsc_douta, din_0_rsc_req_vz, din_0_rsc_rls_lz, din_1_rsc_csa_n, din_1_rsc_csb_n,
      din_1_rsc_addra, din_1_rsc_addrb, din_1_rsc_dinb, din_1_rsc_douta, din_1_rsc_req_vz,
      din_1_rsc_rls_lz, din_2_rsc_csa_n, din_2_rsc_csb_n, din_2_rsc_addra, din_2_rsc_addrb,
      din_2_rsc_dinb, din_2_rsc_douta, din_2_rsc_req_vz, din_2_rsc_rls_lz, din_3_rsc_csa_n,
      din_3_rsc_csb_n, din_3_rsc_addra, din_3_rsc_addrb, din_3_rsc_dinb, din_3_rsc_douta,
      din_3_rsc_req_vz, din_3_rsc_rls_lz, din_4_rsc_csa_n, din_4_rsc_csb_n, din_4_rsc_addra,
      din_4_rsc_addrb, din_4_rsc_dinb, din_4_rsc_douta, din_4_rsc_req_vz, din_4_rsc_rls_lz,
      din_5_rsc_csa_n, din_5_rsc_csb_n, din_5_rsc_addra, din_5_rsc_addrb, din_5_rsc_dinb,
      din_5_rsc_douta, din_5_rsc_req_vz, din_5_rsc_rls_lz, din_6_rsc_csa_n, din_6_rsc_csb_n,
      din_6_rsc_addra, din_6_rsc_addrb, din_6_rsc_dinb, din_6_rsc_douta, din_6_rsc_req_vz,
      din_6_rsc_rls_lz, din_7_rsc_csa_n, din_7_rsc_csb_n, din_7_rsc_addra, din_7_rsc_addrb,
      din_7_rsc_dinb, din_7_rsc_douta, din_7_rsc_req_vz, din_7_rsc_rls_lz, din_8_rsc_csa_n,
      din_8_rsc_csb_n, din_8_rsc_addra, din_8_rsc_addrb, din_8_rsc_dinb, din_8_rsc_douta,
      din_8_rsc_req_vz, din_8_rsc_rls_lz, din_9_rsc_csa_n, din_9_rsc_csb_n, din_9_rsc_addra,
      din_9_rsc_addrb, din_9_rsc_dinb, din_9_rsc_douta, din_9_rsc_req_vz, din_9_rsc_rls_lz,
      din_10_rsc_csa_n, din_10_rsc_csb_n, din_10_rsc_addra, din_10_rsc_addrb, din_10_rsc_dinb,
      din_10_rsc_douta, din_10_rsc_req_vz, din_10_rsc_rls_lz, din_11_rsc_csa_n, din_11_rsc_csb_n,
      din_11_rsc_addra, din_11_rsc_addrb, din_11_rsc_dinb, din_11_rsc_douta, din_11_rsc_req_vz,
      din_11_rsc_rls_lz, din_12_rsc_csa_n, din_12_rsc_csb_n, din_12_rsc_addra, din_12_rsc_addrb,
      din_12_rsc_dinb, din_12_rsc_douta, din_12_rsc_req_vz, din_12_rsc_rls_lz, din_13_rsc_csa_n,
      din_13_rsc_csb_n, din_13_rsc_addra, din_13_rsc_addrb, din_13_rsc_dinb, din_13_rsc_douta,
      din_13_rsc_req_vz, din_13_rsc_rls_lz, din_14_rsc_csa_n, din_14_rsc_csb_n, din_14_rsc_addra,
      din_14_rsc_addrb, din_14_rsc_dinb, din_14_rsc_douta, din_14_rsc_req_vz, din_14_rsc_rls_lz,
      din_15_rsc_csa_n, din_15_rsc_csb_n, din_15_rsc_addra, din_15_rsc_addrb, din_15_rsc_dinb,
      din_15_rsc_douta, din_15_rsc_req_vz, din_15_rsc_rls_lz, din_16_rsc_csa_n, din_16_rsc_csb_n,
      din_16_rsc_addra, din_16_rsc_addrb, din_16_rsc_dinb, din_16_rsc_douta, din_16_rsc_req_vz,
      din_16_rsc_rls_lz, din_17_rsc_csa_n, din_17_rsc_csb_n, din_17_rsc_addra, din_17_rsc_addrb,
      din_17_rsc_dinb, din_17_rsc_douta, din_17_rsc_req_vz, din_17_rsc_rls_lz, dout_rsc_z,
      dout_rsc_vz, dout_rsc_lz
);
  input clk;
  input rst;
  output din_0_rsc_csa_n;
  output din_0_rsc_csb_n;
  output [6:0] din_0_rsc_addra;
  output [6:0] din_0_rsc_addrb;
  output [63:0] din_0_rsc_dinb;
  input [63:0] din_0_rsc_douta;
  input din_0_rsc_req_vz;
  output din_0_rsc_rls_lz;
  output din_1_rsc_csa_n;
  output din_1_rsc_csb_n;
  output [6:0] din_1_rsc_addra;
  output [6:0] din_1_rsc_addrb;
  output [63:0] din_1_rsc_dinb;
  input [63:0] din_1_rsc_douta;
  input din_1_rsc_req_vz;
  output din_1_rsc_rls_lz;
  output din_2_rsc_csa_n;
  output din_2_rsc_csb_n;
  output [6:0] din_2_rsc_addra;
  output [6:0] din_2_rsc_addrb;
  output [63:0] din_2_rsc_dinb;
  input [63:0] din_2_rsc_douta;
  input din_2_rsc_req_vz;
  output din_2_rsc_rls_lz;
  output din_3_rsc_csa_n;
  output din_3_rsc_csb_n;
  output [6:0] din_3_rsc_addra;
  output [6:0] din_3_rsc_addrb;
  output [63:0] din_3_rsc_dinb;
  input [63:0] din_3_rsc_douta;
  input din_3_rsc_req_vz;
  output din_3_rsc_rls_lz;
  output din_4_rsc_csa_n;
  output din_4_rsc_csb_n;
  output [6:0] din_4_rsc_addra;
  output [6:0] din_4_rsc_addrb;
  output [63:0] din_4_rsc_dinb;
  input [63:0] din_4_rsc_douta;
  input din_4_rsc_req_vz;
  output din_4_rsc_rls_lz;
  output din_5_rsc_csa_n;
  output din_5_rsc_csb_n;
  output [6:0] din_5_rsc_addra;
  output [6:0] din_5_rsc_addrb;
  output [63:0] din_5_rsc_dinb;
  input [63:0] din_5_rsc_douta;
  input din_5_rsc_req_vz;
  output din_5_rsc_rls_lz;
  output din_6_rsc_csa_n;
  output din_6_rsc_csb_n;
  output [6:0] din_6_rsc_addra;
  output [6:0] din_6_rsc_addrb;
  output [63:0] din_6_rsc_dinb;
  input [63:0] din_6_rsc_douta;
  input din_6_rsc_req_vz;
  output din_6_rsc_rls_lz;
  output din_7_rsc_csa_n;
  output din_7_rsc_csb_n;
  output [6:0] din_7_rsc_addra;
  output [6:0] din_7_rsc_addrb;
  output [63:0] din_7_rsc_dinb;
  input [63:0] din_7_rsc_douta;
  input din_7_rsc_req_vz;
  output din_7_rsc_rls_lz;
  output din_8_rsc_csa_n;
  output din_8_rsc_csb_n;
  output [6:0] din_8_rsc_addra;
  output [6:0] din_8_rsc_addrb;
  output [63:0] din_8_rsc_dinb;
  input [63:0] din_8_rsc_douta;
  input din_8_rsc_req_vz;
  output din_8_rsc_rls_lz;
  output din_9_rsc_csa_n;
  output din_9_rsc_csb_n;
  output [6:0] din_9_rsc_addra;
  output [6:0] din_9_rsc_addrb;
  output [63:0] din_9_rsc_dinb;
  input [63:0] din_9_rsc_douta;
  input din_9_rsc_req_vz;
  output din_9_rsc_rls_lz;
  output din_10_rsc_csa_n;
  output din_10_rsc_csb_n;
  output [6:0] din_10_rsc_addra;
  output [6:0] din_10_rsc_addrb;
  output [63:0] din_10_rsc_dinb;
  input [63:0] din_10_rsc_douta;
  input din_10_rsc_req_vz;
  output din_10_rsc_rls_lz;
  output din_11_rsc_csa_n;
  output din_11_rsc_csb_n;
  output [6:0] din_11_rsc_addra;
  output [6:0] din_11_rsc_addrb;
  output [63:0] din_11_rsc_dinb;
  input [63:0] din_11_rsc_douta;
  input din_11_rsc_req_vz;
  output din_11_rsc_rls_lz;
  output din_12_rsc_csa_n;
  output din_12_rsc_csb_n;
  output [6:0] din_12_rsc_addra;
  output [6:0] din_12_rsc_addrb;
  output [63:0] din_12_rsc_dinb;
  input [63:0] din_12_rsc_douta;
  input din_12_rsc_req_vz;
  output din_12_rsc_rls_lz;
  output din_13_rsc_csa_n;
  output din_13_rsc_csb_n;
  output [6:0] din_13_rsc_addra;
  output [6:0] din_13_rsc_addrb;
  output [63:0] din_13_rsc_dinb;
  input [63:0] din_13_rsc_douta;
  input din_13_rsc_req_vz;
  output din_13_rsc_rls_lz;
  output din_14_rsc_csa_n;
  output din_14_rsc_csb_n;
  output [6:0] din_14_rsc_addra;
  output [6:0] din_14_rsc_addrb;
  output [63:0] din_14_rsc_dinb;
  input [63:0] din_14_rsc_douta;
  input din_14_rsc_req_vz;
  output din_14_rsc_rls_lz;
  output din_15_rsc_csa_n;
  output din_15_rsc_csb_n;
  output [6:0] din_15_rsc_addra;
  output [6:0] din_15_rsc_addrb;
  output [63:0] din_15_rsc_dinb;
  input [63:0] din_15_rsc_douta;
  input din_15_rsc_req_vz;
  output din_15_rsc_rls_lz;
  output din_16_rsc_csa_n;
  output din_16_rsc_csb_n;
  output [6:0] din_16_rsc_addra;
  output [6:0] din_16_rsc_addrb;
  output [63:0] din_16_rsc_dinb;
  input [63:0] din_16_rsc_douta;
  input din_16_rsc_req_vz;
  output din_16_rsc_rls_lz;
  output din_17_rsc_csa_n;
  output din_17_rsc_csb_n;
  output [6:0] din_17_rsc_addra;
  output [6:0] din_17_rsc_addrb;
  output [63:0] din_17_rsc_dinb;
  input [63:0] din_17_rsc_douta;
  input din_17_rsc_req_vz;
  output din_17_rsc_rls_lz;
  output [511:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;


  // Interconnect Declarations
  wire [63:0] din_0_rsci_douta_d;
  wire din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_1_rsci_douta_d;
  wire din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_2_rsci_douta_d;
  wire din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_3_rsci_douta_d;
  wire din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_4_rsci_douta_d;
  wire din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_5_rsci_douta_d;
  wire din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_6_rsci_douta_d;
  wire din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_7_rsci_douta_d;
  wire din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_8_rsci_douta_d;
  wire din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_9_rsci_douta_d;
  wire din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_10_rsci_douta_d;
  wire din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_11_rsci_douta_d;
  wire din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_12_rsci_douta_d;
  wire din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_13_rsci_douta_d;
  wire din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_14_rsci_douta_d;
  wire din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_15_rsci_douta_d;
  wire din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_16_rsci_douta_d;
  wire din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] din_17_rsci_douta_d;
  wire din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [6:0] din_0_rsci_addra_d_iff;


  // Interconnect Declarations for Component Instantiations 
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_38_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_0_rsci (
      .douta(din_0_rsc_douta),
      .dinb(din_0_rsc_dinb),
      .addrb(din_0_rsc_addrb),
      .addra(din_0_rsc_addra),
      .csb_n(din_0_rsc_csb_n),
      .csa_n(din_0_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_0_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_39_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_1_rsci (
      .douta(din_1_rsc_douta),
      .dinb(din_1_rsc_dinb),
      .addrb(din_1_rsc_addrb),
      .addra(din_1_rsc_addra),
      .csb_n(din_1_rsc_csb_n),
      .csa_n(din_1_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_1_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_40_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_2_rsci (
      .douta(din_2_rsc_douta),
      .dinb(din_2_rsc_dinb),
      .addrb(din_2_rsc_addrb),
      .addra(din_2_rsc_addra),
      .csb_n(din_2_rsc_csb_n),
      .csa_n(din_2_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_2_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_41_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_3_rsci (
      .douta(din_3_rsc_douta),
      .dinb(din_3_rsc_dinb),
      .addrb(din_3_rsc_addrb),
      .addra(din_3_rsc_addra),
      .csb_n(din_3_rsc_csb_n),
      .csa_n(din_3_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_3_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_42_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_4_rsci (
      .douta(din_4_rsc_douta),
      .dinb(din_4_rsc_dinb),
      .addrb(din_4_rsc_addrb),
      .addra(din_4_rsc_addra),
      .csb_n(din_4_rsc_csb_n),
      .csa_n(din_4_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_4_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_43_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_5_rsci (
      .douta(din_5_rsc_douta),
      .dinb(din_5_rsc_dinb),
      .addrb(din_5_rsc_addrb),
      .addra(din_5_rsc_addra),
      .csb_n(din_5_rsc_csb_n),
      .csa_n(din_5_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_5_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_44_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_6_rsci (
      .douta(din_6_rsc_douta),
      .dinb(din_6_rsc_dinb),
      .addrb(din_6_rsc_addrb),
      .addra(din_6_rsc_addra),
      .csb_n(din_6_rsc_csb_n),
      .csa_n(din_6_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_6_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_45_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_7_rsci (
      .douta(din_7_rsc_douta),
      .dinb(din_7_rsc_dinb),
      .addrb(din_7_rsc_addrb),
      .addra(din_7_rsc_addra),
      .csb_n(din_7_rsc_csb_n),
      .csa_n(din_7_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_7_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_46_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_8_rsci (
      .douta(din_8_rsc_douta),
      .dinb(din_8_rsc_dinb),
      .addrb(din_8_rsc_addrb),
      .addra(din_8_rsc_addra),
      .csb_n(din_8_rsc_csb_n),
      .csa_n(din_8_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_8_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_47_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_9_rsci (
      .douta(din_9_rsc_douta),
      .dinb(din_9_rsc_dinb),
      .addrb(din_9_rsc_addrb),
      .addra(din_9_rsc_addra),
      .csb_n(din_9_rsc_csb_n),
      .csa_n(din_9_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_9_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_48_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_10_rsci (
      .douta(din_10_rsc_douta),
      .dinb(din_10_rsc_dinb),
      .addrb(din_10_rsc_addrb),
      .addra(din_10_rsc_addra),
      .csb_n(din_10_rsc_csb_n),
      .csa_n(din_10_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_10_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_49_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_11_rsci (
      .douta(din_11_rsc_douta),
      .dinb(din_11_rsc_dinb),
      .addrb(din_11_rsc_addrb),
      .addra(din_11_rsc_addra),
      .csb_n(din_11_rsc_csb_n),
      .csa_n(din_11_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_11_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_50_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_12_rsci (
      .douta(din_12_rsc_douta),
      .dinb(din_12_rsc_dinb),
      .addrb(din_12_rsc_addrb),
      .addra(din_12_rsc_addra),
      .csb_n(din_12_rsc_csb_n),
      .csa_n(din_12_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_12_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_51_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_13_rsci (
      .douta(din_13_rsc_douta),
      .dinb(din_13_rsc_dinb),
      .addrb(din_13_rsc_addrb),
      .addra(din_13_rsc_addra),
      .csb_n(din_13_rsc_csb_n),
      .csa_n(din_13_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_13_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_52_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_14_rsci (
      .douta(din_14_rsc_douta),
      .dinb(din_14_rsc_dinb),
      .addrb(din_14_rsc_addrb),
      .addra(din_14_rsc_addra),
      .csb_n(din_14_rsc_csb_n),
      .csa_n(din_14_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_14_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_53_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_15_rsci (
      .douta(din_15_rsc_douta),
      .dinb(din_15_rsc_dinb),
      .addrb(din_15_rsc_addrb),
      .addra(din_15_rsc_addra),
      .csb_n(din_15_rsc_csb_n),
      .csa_n(din_15_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_15_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_54_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_16_rsci (
      .douta(din_16_rsc_douta),
      .dinb(din_16_rsc_dinb),
      .addrb(din_16_rsc_addrb),
      .addra(din_16_rsc_addra),
      .csb_n(din_16_rsc_csb_n),
      .csa_n(din_16_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_16_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_55_n1073741823_0_0_0_66_16_66_0_0_0_0_0_0_gen
      din_17_rsci (
      .douta(din_17_rsc_douta),
      .dinb(din_17_rsc_dinb),
      .addrb(din_17_rsc_addrb),
      .addra(din_17_rsc_addra),
      .csb_n(din_17_rsc_csb_n),
      .csa_n(din_17_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d_iff),
      .addrb_d(din_0_rsci_addra_d_iff),
      .dinb_d(64'b0),
      .douta_d(din_17_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_core_inst
      (
      .clk(clk),
      .rst(rst),
      .din_0_rsc_req_vz(din_0_rsc_req_vz),
      .din_0_rsc_rls_lz(din_0_rsc_rls_lz),
      .din_1_rsc_req_vz(din_1_rsc_req_vz),
      .din_1_rsc_rls_lz(din_1_rsc_rls_lz),
      .din_2_rsc_req_vz(din_2_rsc_req_vz),
      .din_2_rsc_rls_lz(din_2_rsc_rls_lz),
      .din_3_rsc_req_vz(din_3_rsc_req_vz),
      .din_3_rsc_rls_lz(din_3_rsc_rls_lz),
      .din_4_rsc_req_vz(din_4_rsc_req_vz),
      .din_4_rsc_rls_lz(din_4_rsc_rls_lz),
      .din_5_rsc_req_vz(din_5_rsc_req_vz),
      .din_5_rsc_rls_lz(din_5_rsc_rls_lz),
      .din_6_rsc_req_vz(din_6_rsc_req_vz),
      .din_6_rsc_rls_lz(din_6_rsc_rls_lz),
      .din_7_rsc_req_vz(din_7_rsc_req_vz),
      .din_7_rsc_rls_lz(din_7_rsc_rls_lz),
      .din_8_rsc_req_vz(din_8_rsc_req_vz),
      .din_8_rsc_rls_lz(din_8_rsc_rls_lz),
      .din_9_rsc_req_vz(din_9_rsc_req_vz),
      .din_9_rsc_rls_lz(din_9_rsc_rls_lz),
      .din_10_rsc_req_vz(din_10_rsc_req_vz),
      .din_10_rsc_rls_lz(din_10_rsc_rls_lz),
      .din_11_rsc_req_vz(din_11_rsc_req_vz),
      .din_11_rsc_rls_lz(din_11_rsc_rls_lz),
      .din_12_rsc_req_vz(din_12_rsc_req_vz),
      .din_12_rsc_rls_lz(din_12_rsc_rls_lz),
      .din_13_rsc_req_vz(din_13_rsc_req_vz),
      .din_13_rsc_rls_lz(din_13_rsc_rls_lz),
      .din_14_rsc_req_vz(din_14_rsc_req_vz),
      .din_14_rsc_rls_lz(din_14_rsc_rls_lz),
      .din_15_rsc_req_vz(din_15_rsc_req_vz),
      .din_15_rsc_rls_lz(din_15_rsc_rls_lz),
      .din_16_rsc_req_vz(din_16_rsc_req_vz),
      .din_16_rsc_rls_lz(din_16_rsc_rls_lz),
      .din_17_rsc_req_vz(din_17_rsc_req_vz),
      .din_17_rsc_rls_lz(din_17_rsc_rls_lz),
      .dout_rsc_z(dout_rsc_z),
      .dout_rsc_vz(dout_rsc_vz),
      .dout_rsc_lz(dout_rsc_lz),
      .din_0_rsci_douta_d(din_0_rsci_douta_d),
      .din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_1_rsci_douta_d(din_1_rsci_douta_d),
      .din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_2_rsci_douta_d(din_2_rsci_douta_d),
      .din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_3_rsci_douta_d(din_3_rsci_douta_d),
      .din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_4_rsci_douta_d(din_4_rsci_douta_d),
      .din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_5_rsci_douta_d(din_5_rsci_douta_d),
      .din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_6_rsci_douta_d(din_6_rsci_douta_d),
      .din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_7_rsci_douta_d(din_7_rsci_douta_d),
      .din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_8_rsci_douta_d(din_8_rsci_douta_d),
      .din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_9_rsci_douta_d(din_9_rsci_douta_d),
      .din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_10_rsci_douta_d(din_10_rsci_douta_d),
      .din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_11_rsci_douta_d(din_11_rsci_douta_d),
      .din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_12_rsci_douta_d(din_12_rsci_douta_d),
      .din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_13_rsci_douta_d(din_13_rsci_douta_d),
      .din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_14_rsci_douta_d(din_14_rsci_douta_d),
      .din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_15_rsci_douta_d(din_15_rsci_douta_d),
      .din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_16_rsci_douta_d(din_16_rsci_douta_d),
      .din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_16_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_17_rsci_douta_d(din_17_rsci_douta_d),
      .din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_17_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_0_rsci_addra_d_pff(din_0_rsci_addra_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_1
// ------------------------------------------------------------------


module WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_1 (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, dout_rsc_csa_n, dout_rsc_csb_n, dout_rsc_addra,
      dout_rsc_addrb, dout_rsc_dinb, dout_rsc_douta, dout_rsc_req_vz, dout_rsc_rls_lz
);
  input clk;
  input rst;
  input [63:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  output dout_rsc_csa_n;
  output dout_rsc_csb_n;
  output [6:0] dout_rsc_addra;
  output [6:0] dout_rsc_addrb;
  output [63:0] dout_rsc_dinb;
  input [63:0] dout_rsc_douta;
  input dout_rsc_req_vz;
  output dout_rsc_rls_lz;


  // Interconnect Declarations
  wire [6:0] dout_rsci_addra_d;
  wire [6:0] dout_rsci_addrb_d;
  wire [63:0] dout_rsci_dinb_d;
  wire [63:0] dout_rsci_douta_d;
  wire dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_96_n1073741823_0_0_0_36_64_128_0_0_0_0_0_0_gen
      dout_rsci (
      .douta(dout_rsc_douta),
      .dinb(dout_rsc_dinb),
      .addrb(dout_rsc_addrb),
      .addra(dout_rsc_addra),
      .csb_n(dout_rsc_csb_n),
      .csa_n(dout_rsc_csa_n),
      .addra_d(dout_rsci_addra_d),
      .addrb_d(dout_rsci_addrb_d),
      .dinb_d(dout_rsci_dinb_d),
      .douta_d(dout_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_core_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(din_rsc_z),
      .din_rsc_vz(din_rsc_vz),
      .din_rsc_lz(din_rsc_lz),
      .dout_rsc_req_vz(dout_rsc_req_vz),
      .dout_rsc_rls_lz(dout_rsc_rls_lz),
      .dout_rsci_addra_d(dout_rsci_addra_d),
      .dout_rsci_addrb_d(dout_rsci_addrb_d),
      .dout_rsci_dinb_d(dout_rsci_dinb_d),
      .dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_1
// ------------------------------------------------------------------


module READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_1 (
  clk, rst, din_rsc_csa_n, din_rsc_csb_n, din_rsc_addra, din_rsc_addrb, din_rsc_dinb,
      din_rsc_douta, din_rsc_req_vz, din_rsc_rls_lz, dout_rsc_z, dout_rsc_vz, dout_rsc_lz
);
  input clk;
  input rst;
  output din_rsc_csa_n;
  output din_rsc_csb_n;
  output [6:0] din_rsc_addra;
  output [6:0] din_rsc_addrb;
  output [63:0] din_rsc_dinb;
  input [63:0] din_rsc_douta;
  input din_rsc_req_vz;
  output din_rsc_rls_lz;
  output [63:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;


  // Interconnect Declarations
  wire [6:0] din_rsci_addra_d;
  wire [6:0] din_rsci_addrb_d;
  wire [63:0] din_rsci_douta_d;
  wire din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  catapult_2p_half_memory_128x64_065nm_cat_ram2p_half_128x64_rwport_98_n1073741823_0_0_0_36_64_128_0_0_0_0_0_0_gen
      din_rsci (
      .douta(din_rsc_douta),
      .dinb(din_rsc_dinb),
      .addrb(din_rsc_addrb),
      .addra(din_rsc_addra),
      .csb_n(din_rsc_csb_n),
      .csa_n(din_rsc_csa_n),
      .addra_d(din_rsci_addra_d),
      .addrb_d(din_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_core_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_req_vz(din_rsc_req_vz),
      .din_rsc_rls_lz(din_rsc_rls_lz),
      .dout_rsc_z(dout_rsc_z),
      .dout_rsc_vz(dout_rsc_vz),
      .dout_rsc_lz(dout_rsc_lz),
      .din_rsci_addra_d(din_rsci_addra_d),
      .din_rsci_addrb_d(din_rsci_addrb_d),
      .din_rsci_douta_d(din_rsci_douta_d),
      .din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    systolic_array
// ------------------------------------------------------------------


module systolic_array (
  clk, rst, input_rsc_z, input_rsc_vz, input_rsc_lz, weight_rsc_z, weight_rsc_vz,
      weight_rsc_lz, output_rsc_z, output_rsc_vz, output_rsc_lz
);
  input clk;
  input rst;
  input [511:0] input_rsc_z;
  input input_rsc_vz;
  output input_rsc_lz;
  input [63:0] weight_rsc_z;
  input weight_rsc_vz;
  output weight_rsc_lz;
  output [1023:0] output_rsc_z;
  input output_rsc_vz;
  output output_rsc_lz;



  // Interconnect Declarations for Component Instantiations 
  systolic_array_core systolic_array_core_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_z(input_rsc_z),
      .input_rsc_vz(input_rsc_vz),
      .input_rsc_lz(input_rsc_lz),
      .weight_rsc_z(weight_rsc_z),
      .weight_rsc_vz(weight_rsc_vz),
      .weight_rsc_lz(weight_rsc_lz),
      .output_rsc_z(output_rsc_z),
      .output_rsc_vz(output_rsc_vz),
      .output_rsc_lz(output_rsc_lz)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_1
// ------------------------------------------------------------------


module WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_1 (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, dout_0_rsc_csa_n, dout_0_rsc_csb_n,
      dout_0_rsc_addra, dout_0_rsc_addrb, dout_0_rsc_dinb, dout_0_rsc_douta, dout_0_rsc_req_vz,
      dout_0_rsc_rls_lz, dout_1_rsc_csa_n, dout_1_rsc_csb_n, dout_1_rsc_addra, dout_1_rsc_addrb,
      dout_1_rsc_dinb, dout_1_rsc_douta, dout_1_rsc_req_vz, dout_1_rsc_rls_lz, dout_2_rsc_csa_n,
      dout_2_rsc_csb_n, dout_2_rsc_addra, dout_2_rsc_addrb, dout_2_rsc_dinb, dout_2_rsc_douta,
      dout_2_rsc_req_vz, dout_2_rsc_rls_lz, dout_3_rsc_csa_n, dout_3_rsc_csb_n, dout_3_rsc_addra,
      dout_3_rsc_addrb, dout_3_rsc_dinb, dout_3_rsc_douta, dout_3_rsc_req_vz, dout_3_rsc_rls_lz,
      dout_4_rsc_csa_n, dout_4_rsc_csb_n, dout_4_rsc_addra, dout_4_rsc_addrb, dout_4_rsc_dinb,
      dout_4_rsc_douta, dout_4_rsc_req_vz, dout_4_rsc_rls_lz, dout_5_rsc_csa_n, dout_5_rsc_csb_n,
      dout_5_rsc_addra, dout_5_rsc_addrb, dout_5_rsc_dinb, dout_5_rsc_douta, dout_5_rsc_req_vz,
      dout_5_rsc_rls_lz, dout_6_rsc_csa_n, dout_6_rsc_csb_n, dout_6_rsc_addra, dout_6_rsc_addrb,
      dout_6_rsc_dinb, dout_6_rsc_douta, dout_6_rsc_req_vz, dout_6_rsc_rls_lz, dout_7_rsc_csa_n,
      dout_7_rsc_csb_n, dout_7_rsc_addra, dout_7_rsc_addrb, dout_7_rsc_dinb, dout_7_rsc_douta,
      dout_7_rsc_req_vz, dout_7_rsc_rls_lz, dout_8_rsc_csa_n, dout_8_rsc_csb_n, dout_8_rsc_addra,
      dout_8_rsc_addrb, dout_8_rsc_dinb, dout_8_rsc_douta, dout_8_rsc_req_vz, dout_8_rsc_rls_lz,
      dout_9_rsc_csa_n, dout_9_rsc_csb_n, dout_9_rsc_addra, dout_9_rsc_addrb, dout_9_rsc_dinb,
      dout_9_rsc_douta, dout_9_rsc_req_vz, dout_9_rsc_rls_lz, dout_10_rsc_csa_n,
      dout_10_rsc_csb_n, dout_10_rsc_addra, dout_10_rsc_addrb, dout_10_rsc_dinb,
      dout_10_rsc_douta, dout_10_rsc_req_vz, dout_10_rsc_rls_lz, dout_11_rsc_csa_n,
      dout_11_rsc_csb_n, dout_11_rsc_addra, dout_11_rsc_addrb, dout_11_rsc_dinb,
      dout_11_rsc_douta, dout_11_rsc_req_vz, dout_11_rsc_rls_lz, dout_12_rsc_csa_n,
      dout_12_rsc_csb_n, dout_12_rsc_addra, dout_12_rsc_addrb, dout_12_rsc_dinb,
      dout_12_rsc_douta, dout_12_rsc_req_vz, dout_12_rsc_rls_lz, dout_13_rsc_csa_n,
      dout_13_rsc_csb_n, dout_13_rsc_addra, dout_13_rsc_addrb, dout_13_rsc_dinb,
      dout_13_rsc_douta, dout_13_rsc_req_vz, dout_13_rsc_rls_lz, dout_14_rsc_csa_n,
      dout_14_rsc_csb_n, dout_14_rsc_addra, dout_14_rsc_addrb, dout_14_rsc_dinb,
      dout_14_rsc_douta, dout_14_rsc_req_vz, dout_14_rsc_rls_lz, dout_15_rsc_csa_n,
      dout_15_rsc_csb_n, dout_15_rsc_addra, dout_15_rsc_addrb, dout_15_rsc_dinb,
      dout_15_rsc_douta, dout_15_rsc_req_vz, dout_15_rsc_rls_lz
);
  input clk;
  input rst;
  input [1023:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  output dout_0_rsc_csa_n;
  output dout_0_rsc_csb_n;
  output [7:0] dout_0_rsc_addra;
  output [7:0] dout_0_rsc_addrb;
  output [63:0] dout_0_rsc_dinb;
  input [63:0] dout_0_rsc_douta;
  input dout_0_rsc_req_vz;
  output dout_0_rsc_rls_lz;
  output dout_1_rsc_csa_n;
  output dout_1_rsc_csb_n;
  output [7:0] dout_1_rsc_addra;
  output [7:0] dout_1_rsc_addrb;
  output [63:0] dout_1_rsc_dinb;
  input [63:0] dout_1_rsc_douta;
  input dout_1_rsc_req_vz;
  output dout_1_rsc_rls_lz;
  output dout_2_rsc_csa_n;
  output dout_2_rsc_csb_n;
  output [7:0] dout_2_rsc_addra;
  output [7:0] dout_2_rsc_addrb;
  output [63:0] dout_2_rsc_dinb;
  input [63:0] dout_2_rsc_douta;
  input dout_2_rsc_req_vz;
  output dout_2_rsc_rls_lz;
  output dout_3_rsc_csa_n;
  output dout_3_rsc_csb_n;
  output [7:0] dout_3_rsc_addra;
  output [7:0] dout_3_rsc_addrb;
  output [63:0] dout_3_rsc_dinb;
  input [63:0] dout_3_rsc_douta;
  input dout_3_rsc_req_vz;
  output dout_3_rsc_rls_lz;
  output dout_4_rsc_csa_n;
  output dout_4_rsc_csb_n;
  output [7:0] dout_4_rsc_addra;
  output [7:0] dout_4_rsc_addrb;
  output [63:0] dout_4_rsc_dinb;
  input [63:0] dout_4_rsc_douta;
  input dout_4_rsc_req_vz;
  output dout_4_rsc_rls_lz;
  output dout_5_rsc_csa_n;
  output dout_5_rsc_csb_n;
  output [7:0] dout_5_rsc_addra;
  output [7:0] dout_5_rsc_addrb;
  output [63:0] dout_5_rsc_dinb;
  input [63:0] dout_5_rsc_douta;
  input dout_5_rsc_req_vz;
  output dout_5_rsc_rls_lz;
  output dout_6_rsc_csa_n;
  output dout_6_rsc_csb_n;
  output [7:0] dout_6_rsc_addra;
  output [7:0] dout_6_rsc_addrb;
  output [63:0] dout_6_rsc_dinb;
  input [63:0] dout_6_rsc_douta;
  input dout_6_rsc_req_vz;
  output dout_6_rsc_rls_lz;
  output dout_7_rsc_csa_n;
  output dout_7_rsc_csb_n;
  output [7:0] dout_7_rsc_addra;
  output [7:0] dout_7_rsc_addrb;
  output [63:0] dout_7_rsc_dinb;
  input [63:0] dout_7_rsc_douta;
  input dout_7_rsc_req_vz;
  output dout_7_rsc_rls_lz;
  output dout_8_rsc_csa_n;
  output dout_8_rsc_csb_n;
  output [7:0] dout_8_rsc_addra;
  output [7:0] dout_8_rsc_addrb;
  output [63:0] dout_8_rsc_dinb;
  input [63:0] dout_8_rsc_douta;
  input dout_8_rsc_req_vz;
  output dout_8_rsc_rls_lz;
  output dout_9_rsc_csa_n;
  output dout_9_rsc_csb_n;
  output [7:0] dout_9_rsc_addra;
  output [7:0] dout_9_rsc_addrb;
  output [63:0] dout_9_rsc_dinb;
  input [63:0] dout_9_rsc_douta;
  input dout_9_rsc_req_vz;
  output dout_9_rsc_rls_lz;
  output dout_10_rsc_csa_n;
  output dout_10_rsc_csb_n;
  output [7:0] dout_10_rsc_addra;
  output [7:0] dout_10_rsc_addrb;
  output [63:0] dout_10_rsc_dinb;
  input [63:0] dout_10_rsc_douta;
  input dout_10_rsc_req_vz;
  output dout_10_rsc_rls_lz;
  output dout_11_rsc_csa_n;
  output dout_11_rsc_csb_n;
  output [7:0] dout_11_rsc_addra;
  output [7:0] dout_11_rsc_addrb;
  output [63:0] dout_11_rsc_dinb;
  input [63:0] dout_11_rsc_douta;
  input dout_11_rsc_req_vz;
  output dout_11_rsc_rls_lz;
  output dout_12_rsc_csa_n;
  output dout_12_rsc_csb_n;
  output [7:0] dout_12_rsc_addra;
  output [7:0] dout_12_rsc_addrb;
  output [63:0] dout_12_rsc_dinb;
  input [63:0] dout_12_rsc_douta;
  input dout_12_rsc_req_vz;
  output dout_12_rsc_rls_lz;
  output dout_13_rsc_csa_n;
  output dout_13_rsc_csb_n;
  output [7:0] dout_13_rsc_addra;
  output [7:0] dout_13_rsc_addrb;
  output [63:0] dout_13_rsc_dinb;
  input [63:0] dout_13_rsc_douta;
  input dout_13_rsc_req_vz;
  output dout_13_rsc_rls_lz;
  output dout_14_rsc_csa_n;
  output dout_14_rsc_csb_n;
  output [7:0] dout_14_rsc_addra;
  output [7:0] dout_14_rsc_addrb;
  output [63:0] dout_14_rsc_dinb;
  input [63:0] dout_14_rsc_douta;
  input dout_14_rsc_req_vz;
  output dout_14_rsc_rls_lz;
  output dout_15_rsc_csa_n;
  output dout_15_rsc_csb_n;
  output [7:0] dout_15_rsc_addra;
  output [7:0] dout_15_rsc_addrb;
  output [63:0] dout_15_rsc_dinb;
  input [63:0] dout_15_rsc_douta;
  input dout_15_rsc_req_vz;
  output dout_15_rsc_rls_lz;


  // Interconnect Declarations
  wire [7:0] dout_0_rsci_addra_d;
  wire [7:0] dout_0_rsci_addrb_d;
  wire [63:0] dout_0_rsci_dinb_d;
  wire [63:0] dout_0_rsci_douta_d;
  wire dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_1_rsci_addra_d;
  wire [7:0] dout_1_rsci_addrb_d;
  wire [63:0] dout_1_rsci_dinb_d;
  wire [63:0] dout_1_rsci_douta_d;
  wire dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_2_rsci_addra_d;
  wire [7:0] dout_2_rsci_addrb_d;
  wire [63:0] dout_2_rsci_dinb_d;
  wire [63:0] dout_2_rsci_douta_d;
  wire dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_3_rsci_addra_d;
  wire [7:0] dout_3_rsci_addrb_d;
  wire [63:0] dout_3_rsci_dinb_d;
  wire [63:0] dout_3_rsci_douta_d;
  wire dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_4_rsci_addra_d;
  wire [7:0] dout_4_rsci_addrb_d;
  wire [63:0] dout_4_rsci_dinb_d;
  wire [63:0] dout_4_rsci_douta_d;
  wire dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_5_rsci_addra_d;
  wire [7:0] dout_5_rsci_addrb_d;
  wire [63:0] dout_5_rsci_dinb_d;
  wire [63:0] dout_5_rsci_douta_d;
  wire dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_6_rsci_addra_d;
  wire [7:0] dout_6_rsci_addrb_d;
  wire [63:0] dout_6_rsci_dinb_d;
  wire [63:0] dout_6_rsci_douta_d;
  wire dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_7_rsci_addra_d;
  wire [7:0] dout_7_rsci_addrb_d;
  wire [63:0] dout_7_rsci_dinb_d;
  wire [63:0] dout_7_rsci_douta_d;
  wire dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_8_rsci_addra_d;
  wire [7:0] dout_8_rsci_addrb_d;
  wire [63:0] dout_8_rsci_dinb_d;
  wire [63:0] dout_8_rsci_douta_d;
  wire dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_9_rsci_addra_d;
  wire [7:0] dout_9_rsci_addrb_d;
  wire [63:0] dout_9_rsci_dinb_d;
  wire [63:0] dout_9_rsci_douta_d;
  wire dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_10_rsci_addra_d;
  wire [7:0] dout_10_rsci_addrb_d;
  wire [63:0] dout_10_rsci_dinb_d;
  wire [63:0] dout_10_rsci_douta_d;
  wire dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_11_rsci_addra_d;
  wire [7:0] dout_11_rsci_addrb_d;
  wire [63:0] dout_11_rsci_dinb_d;
  wire [63:0] dout_11_rsci_douta_d;
  wire dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_12_rsci_addra_d;
  wire [7:0] dout_12_rsci_addrb_d;
  wire [63:0] dout_12_rsci_dinb_d;
  wire [63:0] dout_12_rsci_douta_d;
  wire dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_13_rsci_addra_d;
  wire [7:0] dout_13_rsci_addrb_d;
  wire [63:0] dout_13_rsci_dinb_d;
  wire [63:0] dout_13_rsci_douta_d;
  wire dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_14_rsci_addra_d;
  wire [7:0] dout_14_rsci_addrb_d;
  wire [63:0] dout_14_rsci_dinb_d;
  wire [63:0] dout_14_rsci_douta_d;
  wire dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [7:0] dout_15_rsci_addra_d;
  wire [7:0] dout_15_rsci_addrb_d;
  wire [63:0] dout_15_rsci_dinb_d;
  wire [63:0] dout_15_rsci_douta_d;
  wire dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_113_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_0_rsci (
      .douta(dout_0_rsc_douta),
      .dinb(dout_0_rsc_dinb),
      .addrb(dout_0_rsc_addrb),
      .addra(dout_0_rsc_addra),
      .csb_n(dout_0_rsc_csb_n),
      .csa_n(dout_0_rsc_csa_n),
      .addra_d(dout_0_rsci_addra_d),
      .addrb_d(dout_0_rsci_addrb_d),
      .dinb_d(dout_0_rsci_dinb_d),
      .douta_d(dout_0_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_114_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_1_rsci (
      .douta(dout_1_rsc_douta),
      .dinb(dout_1_rsc_dinb),
      .addrb(dout_1_rsc_addrb),
      .addra(dout_1_rsc_addra),
      .csb_n(dout_1_rsc_csb_n),
      .csa_n(dout_1_rsc_csa_n),
      .addra_d(dout_1_rsci_addra_d),
      .addrb_d(dout_1_rsci_addrb_d),
      .dinb_d(dout_1_rsci_dinb_d),
      .douta_d(dout_1_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_115_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_2_rsci (
      .douta(dout_2_rsc_douta),
      .dinb(dout_2_rsc_dinb),
      .addrb(dout_2_rsc_addrb),
      .addra(dout_2_rsc_addra),
      .csb_n(dout_2_rsc_csb_n),
      .csa_n(dout_2_rsc_csa_n),
      .addra_d(dout_2_rsci_addra_d),
      .addrb_d(dout_2_rsci_addrb_d),
      .dinb_d(dout_2_rsci_dinb_d),
      .douta_d(dout_2_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_116_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_3_rsci (
      .douta(dout_3_rsc_douta),
      .dinb(dout_3_rsc_dinb),
      .addrb(dout_3_rsc_addrb),
      .addra(dout_3_rsc_addra),
      .csb_n(dout_3_rsc_csb_n),
      .csa_n(dout_3_rsc_csa_n),
      .addra_d(dout_3_rsci_addra_d),
      .addrb_d(dout_3_rsci_addrb_d),
      .dinb_d(dout_3_rsci_dinb_d),
      .douta_d(dout_3_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_117_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_4_rsci (
      .douta(dout_4_rsc_douta),
      .dinb(dout_4_rsc_dinb),
      .addrb(dout_4_rsc_addrb),
      .addra(dout_4_rsc_addra),
      .csb_n(dout_4_rsc_csb_n),
      .csa_n(dout_4_rsc_csa_n),
      .addra_d(dout_4_rsci_addra_d),
      .addrb_d(dout_4_rsci_addrb_d),
      .dinb_d(dout_4_rsci_dinb_d),
      .douta_d(dout_4_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_118_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_5_rsci (
      .douta(dout_5_rsc_douta),
      .dinb(dout_5_rsc_dinb),
      .addrb(dout_5_rsc_addrb),
      .addra(dout_5_rsc_addra),
      .csb_n(dout_5_rsc_csb_n),
      .csa_n(dout_5_rsc_csa_n),
      .addra_d(dout_5_rsci_addra_d),
      .addrb_d(dout_5_rsci_addrb_d),
      .dinb_d(dout_5_rsci_dinb_d),
      .douta_d(dout_5_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_119_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_6_rsci (
      .douta(dout_6_rsc_douta),
      .dinb(dout_6_rsc_dinb),
      .addrb(dout_6_rsc_addrb),
      .addra(dout_6_rsc_addra),
      .csb_n(dout_6_rsc_csb_n),
      .csa_n(dout_6_rsc_csa_n),
      .addra_d(dout_6_rsci_addra_d),
      .addrb_d(dout_6_rsci_addrb_d),
      .dinb_d(dout_6_rsci_dinb_d),
      .douta_d(dout_6_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_120_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_7_rsci (
      .douta(dout_7_rsc_douta),
      .dinb(dout_7_rsc_dinb),
      .addrb(dout_7_rsc_addrb),
      .addra(dout_7_rsc_addra),
      .csb_n(dout_7_rsc_csb_n),
      .csa_n(dout_7_rsc_csa_n),
      .addra_d(dout_7_rsci_addra_d),
      .addrb_d(dout_7_rsci_addrb_d),
      .dinb_d(dout_7_rsci_dinb_d),
      .douta_d(dout_7_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_121_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_8_rsci (
      .douta(dout_8_rsc_douta),
      .dinb(dout_8_rsc_dinb),
      .addrb(dout_8_rsc_addrb),
      .addra(dout_8_rsc_addra),
      .csb_n(dout_8_rsc_csb_n),
      .csa_n(dout_8_rsc_csa_n),
      .addra_d(dout_8_rsci_addra_d),
      .addrb_d(dout_8_rsci_addrb_d),
      .dinb_d(dout_8_rsci_dinb_d),
      .douta_d(dout_8_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_122_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_9_rsci (
      .douta(dout_9_rsc_douta),
      .dinb(dout_9_rsc_dinb),
      .addrb(dout_9_rsc_addrb),
      .addra(dout_9_rsc_addra),
      .csb_n(dout_9_rsc_csb_n),
      .csa_n(dout_9_rsc_csa_n),
      .addra_d(dout_9_rsci_addra_d),
      .addrb_d(dout_9_rsci_addrb_d),
      .dinb_d(dout_9_rsci_dinb_d),
      .douta_d(dout_9_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_123_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_10_rsci (
      .douta(dout_10_rsc_douta),
      .dinb(dout_10_rsc_dinb),
      .addrb(dout_10_rsc_addrb),
      .addra(dout_10_rsc_addra),
      .csb_n(dout_10_rsc_csb_n),
      .csa_n(dout_10_rsc_csa_n),
      .addra_d(dout_10_rsci_addra_d),
      .addrb_d(dout_10_rsci_addrb_d),
      .dinb_d(dout_10_rsci_dinb_d),
      .douta_d(dout_10_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_124_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_11_rsci (
      .douta(dout_11_rsc_douta),
      .dinb(dout_11_rsc_dinb),
      .addrb(dout_11_rsc_addrb),
      .addra(dout_11_rsc_addra),
      .csb_n(dout_11_rsc_csb_n),
      .csa_n(dout_11_rsc_csa_n),
      .addra_d(dout_11_rsci_addra_d),
      .addrb_d(dout_11_rsci_addrb_d),
      .dinb_d(dout_11_rsci_dinb_d),
      .douta_d(dout_11_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_125_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_12_rsci (
      .douta(dout_12_rsc_douta),
      .dinb(dout_12_rsc_dinb),
      .addrb(dout_12_rsc_addrb),
      .addra(dout_12_rsc_addra),
      .csb_n(dout_12_rsc_csb_n),
      .csa_n(dout_12_rsc_csa_n),
      .addra_d(dout_12_rsci_addra_d),
      .addrb_d(dout_12_rsci_addrb_d),
      .dinb_d(dout_12_rsci_dinb_d),
      .douta_d(dout_12_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_126_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_13_rsci (
      .douta(dout_13_rsc_douta),
      .dinb(dout_13_rsc_dinb),
      .addrb(dout_13_rsc_addrb),
      .addra(dout_13_rsc_addra),
      .csb_n(dout_13_rsc_csb_n),
      .csa_n(dout_13_rsc_csa_n),
      .addra_d(dout_13_rsci_addra_d),
      .addrb_d(dout_13_rsci_addrb_d),
      .dinb_d(dout_13_rsci_dinb_d),
      .douta_d(dout_13_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_127_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_14_rsci (
      .douta(dout_14_rsc_douta),
      .dinb(dout_14_rsc_dinb),
      .addrb(dout_14_rsc_addrb),
      .addra(dout_14_rsc_addra),
      .csb_n(dout_14_rsc_csb_n),
      .csa_n(dout_14_rsc_csa_n),
      .addra_d(dout_14_rsci_addra_d),
      .addrb_d(dout_14_rsci_addrb_d),
      .dinb_d(dout_14_rsci_dinb_d),
      .douta_d(dout_14_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_128_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      dout_15_rsci (
      .douta(dout_15_rsc_douta),
      .dinb(dout_15_rsc_dinb),
      .addrb(dout_15_rsc_addrb),
      .addra(dout_15_rsc_addra),
      .csb_n(dout_15_rsc_csb_n),
      .csa_n(dout_15_rsc_csa_n),
      .addra_d(dout_15_rsci_addra_d),
      .addrb_d(dout_15_rsci_addrb_d),
      .dinb_d(dout_15_rsci_dinb_d),
      .douta_d(dout_15_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(din_rsc_z),
      .din_rsc_vz(din_rsc_vz),
      .din_rsc_lz(din_rsc_lz),
      .dout_0_rsc_req_vz(dout_0_rsc_req_vz),
      .dout_0_rsc_rls_lz(dout_0_rsc_rls_lz),
      .dout_1_rsc_req_vz(dout_1_rsc_req_vz),
      .dout_1_rsc_rls_lz(dout_1_rsc_rls_lz),
      .dout_2_rsc_req_vz(dout_2_rsc_req_vz),
      .dout_2_rsc_rls_lz(dout_2_rsc_rls_lz),
      .dout_3_rsc_req_vz(dout_3_rsc_req_vz),
      .dout_3_rsc_rls_lz(dout_3_rsc_rls_lz),
      .dout_4_rsc_req_vz(dout_4_rsc_req_vz),
      .dout_4_rsc_rls_lz(dout_4_rsc_rls_lz),
      .dout_5_rsc_req_vz(dout_5_rsc_req_vz),
      .dout_5_rsc_rls_lz(dout_5_rsc_rls_lz),
      .dout_6_rsc_req_vz(dout_6_rsc_req_vz),
      .dout_6_rsc_rls_lz(dout_6_rsc_rls_lz),
      .dout_7_rsc_req_vz(dout_7_rsc_req_vz),
      .dout_7_rsc_rls_lz(dout_7_rsc_rls_lz),
      .dout_8_rsc_req_vz(dout_8_rsc_req_vz),
      .dout_8_rsc_rls_lz(dout_8_rsc_rls_lz),
      .dout_9_rsc_req_vz(dout_9_rsc_req_vz),
      .dout_9_rsc_rls_lz(dout_9_rsc_rls_lz),
      .dout_10_rsc_req_vz(dout_10_rsc_req_vz),
      .dout_10_rsc_rls_lz(dout_10_rsc_rls_lz),
      .dout_11_rsc_req_vz(dout_11_rsc_req_vz),
      .dout_11_rsc_rls_lz(dout_11_rsc_rls_lz),
      .dout_12_rsc_req_vz(dout_12_rsc_req_vz),
      .dout_12_rsc_rls_lz(dout_12_rsc_rls_lz),
      .dout_13_rsc_req_vz(dout_13_rsc_req_vz),
      .dout_13_rsc_rls_lz(dout_13_rsc_rls_lz),
      .dout_14_rsc_req_vz(dout_14_rsc_req_vz),
      .dout_14_rsc_rls_lz(dout_14_rsc_rls_lz),
      .dout_15_rsc_req_vz(dout_15_rsc_req_vz),
      .dout_15_rsc_rls_lz(dout_15_rsc_rls_lz),
      .dout_0_rsci_addra_d(dout_0_rsci_addra_d),
      .dout_0_rsci_addrb_d(dout_0_rsci_addrb_d),
      .dout_0_rsci_dinb_d(dout_0_rsci_dinb_d),
      .dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_0_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_1_rsci_addra_d(dout_1_rsci_addra_d),
      .dout_1_rsci_addrb_d(dout_1_rsci_addrb_d),
      .dout_1_rsci_dinb_d(dout_1_rsci_dinb_d),
      .dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_1_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_2_rsci_addra_d(dout_2_rsci_addra_d),
      .dout_2_rsci_addrb_d(dout_2_rsci_addrb_d),
      .dout_2_rsci_dinb_d(dout_2_rsci_dinb_d),
      .dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_2_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_3_rsci_addra_d(dout_3_rsci_addra_d),
      .dout_3_rsci_addrb_d(dout_3_rsci_addrb_d),
      .dout_3_rsci_dinb_d(dout_3_rsci_dinb_d),
      .dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_3_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_4_rsci_addra_d(dout_4_rsci_addra_d),
      .dout_4_rsci_addrb_d(dout_4_rsci_addrb_d),
      .dout_4_rsci_dinb_d(dout_4_rsci_dinb_d),
      .dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_4_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_5_rsci_addra_d(dout_5_rsci_addra_d),
      .dout_5_rsci_addrb_d(dout_5_rsci_addrb_d),
      .dout_5_rsci_dinb_d(dout_5_rsci_dinb_d),
      .dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_5_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_6_rsci_addra_d(dout_6_rsci_addra_d),
      .dout_6_rsci_addrb_d(dout_6_rsci_addrb_d),
      .dout_6_rsci_dinb_d(dout_6_rsci_dinb_d),
      .dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_6_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_7_rsci_addra_d(dout_7_rsci_addra_d),
      .dout_7_rsci_addrb_d(dout_7_rsci_addrb_d),
      .dout_7_rsci_dinb_d(dout_7_rsci_dinb_d),
      .dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_7_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_8_rsci_addra_d(dout_8_rsci_addra_d),
      .dout_8_rsci_addrb_d(dout_8_rsci_addrb_d),
      .dout_8_rsci_dinb_d(dout_8_rsci_dinb_d),
      .dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_8_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_9_rsci_addra_d(dout_9_rsci_addra_d),
      .dout_9_rsci_addrb_d(dout_9_rsci_addrb_d),
      .dout_9_rsci_dinb_d(dout_9_rsci_dinb_d),
      .dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_9_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_10_rsci_addra_d(dout_10_rsci_addra_d),
      .dout_10_rsci_addrb_d(dout_10_rsci_addrb_d),
      .dout_10_rsci_dinb_d(dout_10_rsci_dinb_d),
      .dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_10_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_11_rsci_addra_d(dout_11_rsci_addra_d),
      .dout_11_rsci_addrb_d(dout_11_rsci_addrb_d),
      .dout_11_rsci_dinb_d(dout_11_rsci_dinb_d),
      .dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_11_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_12_rsci_addra_d(dout_12_rsci_addra_d),
      .dout_12_rsci_addrb_d(dout_12_rsci_addrb_d),
      .dout_12_rsci_dinb_d(dout_12_rsci_dinb_d),
      .dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_12_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_13_rsci_addra_d(dout_13_rsci_addra_d),
      .dout_13_rsci_addrb_d(dout_13_rsci_addrb_d),
      .dout_13_rsci_dinb_d(dout_13_rsci_dinb_d),
      .dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_13_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_14_rsci_addra_d(dout_14_rsci_addra_d),
      .dout_14_rsci_addrb_d(dout_14_rsci_addrb_d),
      .dout_14_rsci_dinb_d(dout_14_rsci_dinb_d),
      .dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_14_rsci_port_0_rw_ram_ir_internal_WMASK_B_d),
      .dout_15_rsci_addra_d(dout_15_rsci_addra_d),
      .dout_15_rsci_addrb_d(dout_15_rsci_addrb_d),
      .dout_15_rsci_dinb_d(dout_15_rsci_dinb_d),
      .dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d(dout_15_rsci_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_1
// ------------------------------------------------------------------


module READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_1 (
  clk, rst, din_0_rsc_csa_n, din_0_rsc_csb_n, din_0_rsc_addra, din_0_rsc_addrb, din_0_rsc_dinb,
      din_0_rsc_douta, din_0_rsc_req_vz, din_0_rsc_rls_lz, din_1_rsc_csa_n, din_1_rsc_csb_n,
      din_1_rsc_addra, din_1_rsc_addrb, din_1_rsc_dinb, din_1_rsc_douta, din_1_rsc_req_vz,
      din_1_rsc_rls_lz, din_2_rsc_csa_n, din_2_rsc_csb_n, din_2_rsc_addra, din_2_rsc_addrb,
      din_2_rsc_dinb, din_2_rsc_douta, din_2_rsc_req_vz, din_2_rsc_rls_lz, din_3_rsc_csa_n,
      din_3_rsc_csb_n, din_3_rsc_addra, din_3_rsc_addrb, din_3_rsc_dinb, din_3_rsc_douta,
      din_3_rsc_req_vz, din_3_rsc_rls_lz, din_4_rsc_csa_n, din_4_rsc_csb_n, din_4_rsc_addra,
      din_4_rsc_addrb, din_4_rsc_dinb, din_4_rsc_douta, din_4_rsc_req_vz, din_4_rsc_rls_lz,
      din_5_rsc_csa_n, din_5_rsc_csb_n, din_5_rsc_addra, din_5_rsc_addrb, din_5_rsc_dinb,
      din_5_rsc_douta, din_5_rsc_req_vz, din_5_rsc_rls_lz, din_6_rsc_csa_n, din_6_rsc_csb_n,
      din_6_rsc_addra, din_6_rsc_addrb, din_6_rsc_dinb, din_6_rsc_douta, din_6_rsc_req_vz,
      din_6_rsc_rls_lz, din_7_rsc_csa_n, din_7_rsc_csb_n, din_7_rsc_addra, din_7_rsc_addrb,
      din_7_rsc_dinb, din_7_rsc_douta, din_7_rsc_req_vz, din_7_rsc_rls_lz, din_8_rsc_csa_n,
      din_8_rsc_csb_n, din_8_rsc_addra, din_8_rsc_addrb, din_8_rsc_dinb, din_8_rsc_douta,
      din_8_rsc_req_vz, din_8_rsc_rls_lz, din_9_rsc_csa_n, din_9_rsc_csb_n, din_9_rsc_addra,
      din_9_rsc_addrb, din_9_rsc_dinb, din_9_rsc_douta, din_9_rsc_req_vz, din_9_rsc_rls_lz,
      din_10_rsc_csa_n, din_10_rsc_csb_n, din_10_rsc_addra, din_10_rsc_addrb, din_10_rsc_dinb,
      din_10_rsc_douta, din_10_rsc_req_vz, din_10_rsc_rls_lz, din_11_rsc_csa_n, din_11_rsc_csb_n,
      din_11_rsc_addra, din_11_rsc_addrb, din_11_rsc_dinb, din_11_rsc_douta, din_11_rsc_req_vz,
      din_11_rsc_rls_lz, din_12_rsc_csa_n, din_12_rsc_csb_n, din_12_rsc_addra, din_12_rsc_addrb,
      din_12_rsc_dinb, din_12_rsc_douta, din_12_rsc_req_vz, din_12_rsc_rls_lz, din_13_rsc_csa_n,
      din_13_rsc_csb_n, din_13_rsc_addra, din_13_rsc_addrb, din_13_rsc_dinb, din_13_rsc_douta,
      din_13_rsc_req_vz, din_13_rsc_rls_lz, din_14_rsc_csa_n, din_14_rsc_csb_n, din_14_rsc_addra,
      din_14_rsc_addrb, din_14_rsc_dinb, din_14_rsc_douta, din_14_rsc_req_vz, din_14_rsc_rls_lz,
      din_15_rsc_csa_n, din_15_rsc_csb_n, din_15_rsc_addra, din_15_rsc_addrb, din_15_rsc_dinb,
      din_15_rsc_douta, din_15_rsc_req_vz, din_15_rsc_rls_lz, dout_rsc_z, dout_rsc_vz,
      dout_rsc_lz
);
  input clk;
  input rst;
  output din_0_rsc_csa_n;
  output din_0_rsc_csb_n;
  output [7:0] din_0_rsc_addra;
  output [7:0] din_0_rsc_addrb;
  output [63:0] din_0_rsc_dinb;
  input [63:0] din_0_rsc_douta;
  input din_0_rsc_req_vz;
  output din_0_rsc_rls_lz;
  output din_1_rsc_csa_n;
  output din_1_rsc_csb_n;
  output [7:0] din_1_rsc_addra;
  output [7:0] din_1_rsc_addrb;
  output [63:0] din_1_rsc_dinb;
  input [63:0] din_1_rsc_douta;
  input din_1_rsc_req_vz;
  output din_1_rsc_rls_lz;
  output din_2_rsc_csa_n;
  output din_2_rsc_csb_n;
  output [7:0] din_2_rsc_addra;
  output [7:0] din_2_rsc_addrb;
  output [63:0] din_2_rsc_dinb;
  input [63:0] din_2_rsc_douta;
  input din_2_rsc_req_vz;
  output din_2_rsc_rls_lz;
  output din_3_rsc_csa_n;
  output din_3_rsc_csb_n;
  output [7:0] din_3_rsc_addra;
  output [7:0] din_3_rsc_addrb;
  output [63:0] din_3_rsc_dinb;
  input [63:0] din_3_rsc_douta;
  input din_3_rsc_req_vz;
  output din_3_rsc_rls_lz;
  output din_4_rsc_csa_n;
  output din_4_rsc_csb_n;
  output [7:0] din_4_rsc_addra;
  output [7:0] din_4_rsc_addrb;
  output [63:0] din_4_rsc_dinb;
  input [63:0] din_4_rsc_douta;
  input din_4_rsc_req_vz;
  output din_4_rsc_rls_lz;
  output din_5_rsc_csa_n;
  output din_5_rsc_csb_n;
  output [7:0] din_5_rsc_addra;
  output [7:0] din_5_rsc_addrb;
  output [63:0] din_5_rsc_dinb;
  input [63:0] din_5_rsc_douta;
  input din_5_rsc_req_vz;
  output din_5_rsc_rls_lz;
  output din_6_rsc_csa_n;
  output din_6_rsc_csb_n;
  output [7:0] din_6_rsc_addra;
  output [7:0] din_6_rsc_addrb;
  output [63:0] din_6_rsc_dinb;
  input [63:0] din_6_rsc_douta;
  input din_6_rsc_req_vz;
  output din_6_rsc_rls_lz;
  output din_7_rsc_csa_n;
  output din_7_rsc_csb_n;
  output [7:0] din_7_rsc_addra;
  output [7:0] din_7_rsc_addrb;
  output [63:0] din_7_rsc_dinb;
  input [63:0] din_7_rsc_douta;
  input din_7_rsc_req_vz;
  output din_7_rsc_rls_lz;
  output din_8_rsc_csa_n;
  output din_8_rsc_csb_n;
  output [7:0] din_8_rsc_addra;
  output [7:0] din_8_rsc_addrb;
  output [63:0] din_8_rsc_dinb;
  input [63:0] din_8_rsc_douta;
  input din_8_rsc_req_vz;
  output din_8_rsc_rls_lz;
  output din_9_rsc_csa_n;
  output din_9_rsc_csb_n;
  output [7:0] din_9_rsc_addra;
  output [7:0] din_9_rsc_addrb;
  output [63:0] din_9_rsc_dinb;
  input [63:0] din_9_rsc_douta;
  input din_9_rsc_req_vz;
  output din_9_rsc_rls_lz;
  output din_10_rsc_csa_n;
  output din_10_rsc_csb_n;
  output [7:0] din_10_rsc_addra;
  output [7:0] din_10_rsc_addrb;
  output [63:0] din_10_rsc_dinb;
  input [63:0] din_10_rsc_douta;
  input din_10_rsc_req_vz;
  output din_10_rsc_rls_lz;
  output din_11_rsc_csa_n;
  output din_11_rsc_csb_n;
  output [7:0] din_11_rsc_addra;
  output [7:0] din_11_rsc_addrb;
  output [63:0] din_11_rsc_dinb;
  input [63:0] din_11_rsc_douta;
  input din_11_rsc_req_vz;
  output din_11_rsc_rls_lz;
  output din_12_rsc_csa_n;
  output din_12_rsc_csb_n;
  output [7:0] din_12_rsc_addra;
  output [7:0] din_12_rsc_addrb;
  output [63:0] din_12_rsc_dinb;
  input [63:0] din_12_rsc_douta;
  input din_12_rsc_req_vz;
  output din_12_rsc_rls_lz;
  output din_13_rsc_csa_n;
  output din_13_rsc_csb_n;
  output [7:0] din_13_rsc_addra;
  output [7:0] din_13_rsc_addrb;
  output [63:0] din_13_rsc_dinb;
  input [63:0] din_13_rsc_douta;
  input din_13_rsc_req_vz;
  output din_13_rsc_rls_lz;
  output din_14_rsc_csa_n;
  output din_14_rsc_csb_n;
  output [7:0] din_14_rsc_addra;
  output [7:0] din_14_rsc_addrb;
  output [63:0] din_14_rsc_dinb;
  input [63:0] din_14_rsc_douta;
  input din_14_rsc_req_vz;
  output din_14_rsc_rls_lz;
  output din_15_rsc_csa_n;
  output din_15_rsc_csb_n;
  output [7:0] din_15_rsc_addra;
  output [7:0] din_15_rsc_addrb;
  output [63:0] din_15_rsc_dinb;
  input [63:0] din_15_rsc_douta;
  input din_15_rsc_req_vz;
  output din_15_rsc_rls_lz;
  output [1023:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;


  // Interconnect Declarations
  wire [7:0] din_0_rsci_addra_d;
  wire [7:0] din_0_rsci_addrb_d;
  wire [63:0] din_0_rsci_douta_d;
  wire din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_1_rsci_addra_d;
  wire [7:0] din_1_rsci_addrb_d;
  wire [63:0] din_1_rsci_douta_d;
  wire din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_2_rsci_addra_d;
  wire [7:0] din_2_rsci_addrb_d;
  wire [63:0] din_2_rsci_douta_d;
  wire din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_3_rsci_addra_d;
  wire [7:0] din_3_rsci_addrb_d;
  wire [63:0] din_3_rsci_douta_d;
  wire din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_4_rsci_addra_d;
  wire [7:0] din_4_rsci_addrb_d;
  wire [63:0] din_4_rsci_douta_d;
  wire din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_5_rsci_addra_d;
  wire [7:0] din_5_rsci_addrb_d;
  wire [63:0] din_5_rsci_douta_d;
  wire din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_6_rsci_addra_d;
  wire [7:0] din_6_rsci_addrb_d;
  wire [63:0] din_6_rsci_douta_d;
  wire din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_7_rsci_addra_d;
  wire [7:0] din_7_rsci_addrb_d;
  wire [63:0] din_7_rsci_douta_d;
  wire din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_8_rsci_addra_d;
  wire [7:0] din_8_rsci_addrb_d;
  wire [63:0] din_8_rsci_douta_d;
  wire din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_9_rsci_addra_d;
  wire [7:0] din_9_rsci_addrb_d;
  wire [63:0] din_9_rsci_douta_d;
  wire din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_10_rsci_addra_d;
  wire [7:0] din_10_rsci_addrb_d;
  wire [63:0] din_10_rsci_douta_d;
  wire din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_11_rsci_addra_d;
  wire [7:0] din_11_rsci_addrb_d;
  wire [63:0] din_11_rsci_douta_d;
  wire din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_12_rsci_addra_d;
  wire [7:0] din_12_rsci_addrb_d;
  wire [63:0] din_12_rsci_douta_d;
  wire din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_13_rsci_addra_d;
  wire [7:0] din_13_rsci_addrb_d;
  wire [63:0] din_13_rsci_douta_d;
  wire din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_14_rsci_addra_d;
  wire [7:0] din_14_rsci_addrb_d;
  wire [63:0] din_14_rsci_douta_d;
  wire din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] din_15_rsci_addra_d;
  wire [7:0] din_15_rsci_addrb_d;
  wire [63:0] din_15_rsci_douta_d;
  wire din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_145_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_0_rsci (
      .douta(din_0_rsc_douta),
      .dinb(din_0_rsc_dinb),
      .addrb(din_0_rsc_addrb),
      .addra(din_0_rsc_addra),
      .csb_n(din_0_rsc_csb_n),
      .csa_n(din_0_rsc_csa_n),
      .addra_d(din_0_rsci_addra_d),
      .addrb_d(din_0_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_0_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_146_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_1_rsci (
      .douta(din_1_rsc_douta),
      .dinb(din_1_rsc_dinb),
      .addrb(din_1_rsc_addrb),
      .addra(din_1_rsc_addra),
      .csb_n(din_1_rsc_csb_n),
      .csa_n(din_1_rsc_csa_n),
      .addra_d(din_1_rsci_addra_d),
      .addrb_d(din_1_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_1_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_147_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_2_rsci (
      .douta(din_2_rsc_douta),
      .dinb(din_2_rsc_dinb),
      .addrb(din_2_rsc_addrb),
      .addra(din_2_rsc_addra),
      .csb_n(din_2_rsc_csb_n),
      .csa_n(din_2_rsc_csa_n),
      .addra_d(din_2_rsci_addra_d),
      .addrb_d(din_2_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_2_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_148_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_3_rsci (
      .douta(din_3_rsc_douta),
      .dinb(din_3_rsc_dinb),
      .addrb(din_3_rsc_addrb),
      .addra(din_3_rsc_addra),
      .csb_n(din_3_rsc_csb_n),
      .csa_n(din_3_rsc_csa_n),
      .addra_d(din_3_rsci_addra_d),
      .addrb_d(din_3_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_3_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_149_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_4_rsci (
      .douta(din_4_rsc_douta),
      .dinb(din_4_rsc_dinb),
      .addrb(din_4_rsc_addrb),
      .addra(din_4_rsc_addra),
      .csb_n(din_4_rsc_csb_n),
      .csa_n(din_4_rsc_csa_n),
      .addra_d(din_4_rsci_addra_d),
      .addrb_d(din_4_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_4_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_150_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_5_rsci (
      .douta(din_5_rsc_douta),
      .dinb(din_5_rsc_dinb),
      .addrb(din_5_rsc_addrb),
      .addra(din_5_rsc_addra),
      .csb_n(din_5_rsc_csb_n),
      .csa_n(din_5_rsc_csa_n),
      .addra_d(din_5_rsci_addra_d),
      .addrb_d(din_5_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_5_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_151_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_6_rsci (
      .douta(din_6_rsc_douta),
      .dinb(din_6_rsc_dinb),
      .addrb(din_6_rsc_addrb),
      .addra(din_6_rsc_addra),
      .csb_n(din_6_rsc_csb_n),
      .csa_n(din_6_rsc_csa_n),
      .addra_d(din_6_rsci_addra_d),
      .addrb_d(din_6_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_6_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_152_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_7_rsci (
      .douta(din_7_rsc_douta),
      .dinb(din_7_rsc_dinb),
      .addrb(din_7_rsc_addrb),
      .addra(din_7_rsc_addra),
      .csb_n(din_7_rsc_csb_n),
      .csa_n(din_7_rsc_csa_n),
      .addra_d(din_7_rsci_addra_d),
      .addrb_d(din_7_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_7_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_153_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_8_rsci (
      .douta(din_8_rsc_douta),
      .dinb(din_8_rsc_dinb),
      .addrb(din_8_rsc_addrb),
      .addra(din_8_rsc_addra),
      .csb_n(din_8_rsc_csb_n),
      .csa_n(din_8_rsc_csa_n),
      .addra_d(din_8_rsci_addra_d),
      .addrb_d(din_8_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_8_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_154_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_9_rsci (
      .douta(din_9_rsc_douta),
      .dinb(din_9_rsc_dinb),
      .addrb(din_9_rsc_addrb),
      .addra(din_9_rsc_addra),
      .csb_n(din_9_rsc_csb_n),
      .csa_n(din_9_rsc_csa_n),
      .addra_d(din_9_rsci_addra_d),
      .addrb_d(din_9_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_9_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_155_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_10_rsci (
      .douta(din_10_rsc_douta),
      .dinb(din_10_rsc_dinb),
      .addrb(din_10_rsc_addrb),
      .addra(din_10_rsc_addra),
      .csb_n(din_10_rsc_csb_n),
      .csa_n(din_10_rsc_csa_n),
      .addra_d(din_10_rsci_addra_d),
      .addrb_d(din_10_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_10_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_156_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_11_rsci (
      .douta(din_11_rsc_douta),
      .dinb(din_11_rsc_dinb),
      .addrb(din_11_rsc_addrb),
      .addra(din_11_rsc_addra),
      .csb_n(din_11_rsc_csb_n),
      .csa_n(din_11_rsc_csa_n),
      .addra_d(din_11_rsci_addra_d),
      .addrb_d(din_11_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_11_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_157_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_12_rsci (
      .douta(din_12_rsc_douta),
      .dinb(din_12_rsc_dinb),
      .addrb(din_12_rsc_addrb),
      .addra(din_12_rsc_addra),
      .csb_n(din_12_rsc_csb_n),
      .csa_n(din_12_rsc_csa_n),
      .addra_d(din_12_rsci_addra_d),
      .addrb_d(din_12_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_12_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_158_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_13_rsci (
      .douta(din_13_rsc_douta),
      .dinb(din_13_rsc_dinb),
      .addrb(din_13_rsc_addrb),
      .addra(din_13_rsc_addra),
      .csb_n(din_13_rsc_csb_n),
      .csa_n(din_13_rsc_csa_n),
      .addra_d(din_13_rsci_addra_d),
      .addrb_d(din_13_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_13_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_159_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_14_rsci (
      .douta(din_14_rsc_douta),
      .dinb(din_14_rsc_dinb),
      .addrb(din_14_rsc_addrb),
      .addra(din_14_rsc_addra),
      .csb_n(din_14_rsc_csb_n),
      .csa_n(din_14_rsc_csa_n),
      .addra_d(din_14_rsci_addra_d),
      .addrb_d(din_14_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_14_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  catapult_2p_half_memory_065nm_cat_ram2p_half_rwport_160_n1073741823_n1073741823_256_64_256_0_0_0_0_0_0_0_gen
      din_15_rsci (
      .douta(din_15_rsc_douta),
      .dinb(din_15_rsc_dinb),
      .addrb(din_15_rsc_addrb),
      .addra(din_15_rsc_addra),
      .csb_n(din_15_rsc_csb_n),
      .csa_n(din_15_rsc_csa_n),
      .addra_d(din_15_rsci_addra_d),
      .addrb_d(din_15_rsci_addrb_d),
      .dinb_d(64'b0),
      .douta_d(din_15_rsci_douta_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_core_inst
      (
      .clk(clk),
      .rst(rst),
      .din_0_rsc_req_vz(din_0_rsc_req_vz),
      .din_0_rsc_rls_lz(din_0_rsc_rls_lz),
      .din_1_rsc_req_vz(din_1_rsc_req_vz),
      .din_1_rsc_rls_lz(din_1_rsc_rls_lz),
      .din_2_rsc_req_vz(din_2_rsc_req_vz),
      .din_2_rsc_rls_lz(din_2_rsc_rls_lz),
      .din_3_rsc_req_vz(din_3_rsc_req_vz),
      .din_3_rsc_rls_lz(din_3_rsc_rls_lz),
      .din_4_rsc_req_vz(din_4_rsc_req_vz),
      .din_4_rsc_rls_lz(din_4_rsc_rls_lz),
      .din_5_rsc_req_vz(din_5_rsc_req_vz),
      .din_5_rsc_rls_lz(din_5_rsc_rls_lz),
      .din_6_rsc_req_vz(din_6_rsc_req_vz),
      .din_6_rsc_rls_lz(din_6_rsc_rls_lz),
      .din_7_rsc_req_vz(din_7_rsc_req_vz),
      .din_7_rsc_rls_lz(din_7_rsc_rls_lz),
      .din_8_rsc_req_vz(din_8_rsc_req_vz),
      .din_8_rsc_rls_lz(din_8_rsc_rls_lz),
      .din_9_rsc_req_vz(din_9_rsc_req_vz),
      .din_9_rsc_rls_lz(din_9_rsc_rls_lz),
      .din_10_rsc_req_vz(din_10_rsc_req_vz),
      .din_10_rsc_rls_lz(din_10_rsc_rls_lz),
      .din_11_rsc_req_vz(din_11_rsc_req_vz),
      .din_11_rsc_rls_lz(din_11_rsc_rls_lz),
      .din_12_rsc_req_vz(din_12_rsc_req_vz),
      .din_12_rsc_rls_lz(din_12_rsc_rls_lz),
      .din_13_rsc_req_vz(din_13_rsc_req_vz),
      .din_13_rsc_rls_lz(din_13_rsc_rls_lz),
      .din_14_rsc_req_vz(din_14_rsc_req_vz),
      .din_14_rsc_rls_lz(din_14_rsc_rls_lz),
      .din_15_rsc_req_vz(din_15_rsc_req_vz),
      .din_15_rsc_rls_lz(din_15_rsc_rls_lz),
      .dout_rsc_z(dout_rsc_z),
      .dout_rsc_vz(dout_rsc_vz),
      .dout_rsc_lz(dout_rsc_lz),
      .din_0_rsci_addra_d(din_0_rsci_addra_d),
      .din_0_rsci_addrb_d(din_0_rsci_addrb_d),
      .din_0_rsci_douta_d(din_0_rsci_douta_d),
      .din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_0_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_1_rsci_addra_d(din_1_rsci_addra_d),
      .din_1_rsci_addrb_d(din_1_rsci_addrb_d),
      .din_1_rsci_douta_d(din_1_rsci_douta_d),
      .din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_1_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_2_rsci_addra_d(din_2_rsci_addra_d),
      .din_2_rsci_addrb_d(din_2_rsci_addrb_d),
      .din_2_rsci_douta_d(din_2_rsci_douta_d),
      .din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_2_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_3_rsci_addra_d(din_3_rsci_addra_d),
      .din_3_rsci_addrb_d(din_3_rsci_addrb_d),
      .din_3_rsci_douta_d(din_3_rsci_douta_d),
      .din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_3_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_4_rsci_addra_d(din_4_rsci_addra_d),
      .din_4_rsci_addrb_d(din_4_rsci_addrb_d),
      .din_4_rsci_douta_d(din_4_rsci_douta_d),
      .din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_4_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_5_rsci_addra_d(din_5_rsci_addra_d),
      .din_5_rsci_addrb_d(din_5_rsci_addrb_d),
      .din_5_rsci_douta_d(din_5_rsci_douta_d),
      .din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_5_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_6_rsci_addra_d(din_6_rsci_addra_d),
      .din_6_rsci_addrb_d(din_6_rsci_addrb_d),
      .din_6_rsci_douta_d(din_6_rsci_douta_d),
      .din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_6_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_7_rsci_addra_d(din_7_rsci_addra_d),
      .din_7_rsci_addrb_d(din_7_rsci_addrb_d),
      .din_7_rsci_douta_d(din_7_rsci_douta_d),
      .din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_7_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_8_rsci_addra_d(din_8_rsci_addra_d),
      .din_8_rsci_addrb_d(din_8_rsci_addrb_d),
      .din_8_rsci_douta_d(din_8_rsci_douta_d),
      .din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_8_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_9_rsci_addra_d(din_9_rsci_addra_d),
      .din_9_rsci_addrb_d(din_9_rsci_addrb_d),
      .din_9_rsci_douta_d(din_9_rsci_douta_d),
      .din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_9_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_10_rsci_addra_d(din_10_rsci_addra_d),
      .din_10_rsci_addrb_d(din_10_rsci_addrb_d),
      .din_10_rsci_douta_d(din_10_rsci_douta_d),
      .din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_10_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_11_rsci_addra_d(din_11_rsci_addra_d),
      .din_11_rsci_addrb_d(din_11_rsci_addrb_d),
      .din_11_rsci_douta_d(din_11_rsci_douta_d),
      .din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_11_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_12_rsci_addra_d(din_12_rsci_addra_d),
      .din_12_rsci_addrb_d(din_12_rsci_addrb_d),
      .din_12_rsci_douta_d(din_12_rsci_douta_d),
      .din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_12_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_13_rsci_addra_d(din_13_rsci_addra_d),
      .din_13_rsci_addrb_d(din_13_rsci_addrb_d),
      .din_13_rsci_douta_d(din_13_rsci_douta_d),
      .din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_13_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_14_rsci_addra_d(din_14_rsci_addra_d),
      .din_14_rsci_addrb_d(din_14_rsci_addrb_d),
      .din_14_rsci_douta_d(din_14_rsci_douta_d),
      .din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_14_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .din_15_rsci_addra_d(din_15_rsci_addra_d),
      .din_15_rsci_addrb_d(din_15_rsci_addrb_d),
      .din_15_rsci_douta_d(din_15_rsci_douta_d),
      .din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_15_rsci_port_0_rw_ram_ir_internal_RMASK_B_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffer_input_DTYPE_64_16_4_1_3
// ------------------------------------------------------------------


module double_buffer_input_DTYPE_64_16_4_1_3 (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, dout_rsc_z, dout_rsc_vz, dout_rsc_lz,
      clamp_mem, scan_n, shift_n, slp_nret_n, slp_ret_n
);
  input clk;
  input rst;
  input [15:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  output [511:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;
  input clamp_mem;
  input scan_n;
  input shift_n;
  input slp_nret_n;
  input slp_ret_n;


  // Interconnect Declarations
  wire din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_0_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_0_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_0_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_0_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_0_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_0_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_0_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_1_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_1_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_1_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_1_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_1_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_2_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_2_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_2_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_2_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_2_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_3_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_3_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_3_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_3_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_3_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_4_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_4_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_4_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_4_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_4_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_5_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_5_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_5_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_5_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_5_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_6_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_6_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_6_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_6_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_6_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_7_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_7_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_7_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_7_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_7_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_8_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_8_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_8_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_8_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_8_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_9_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_9_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_9_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_9_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_9_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_10_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_10_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_10_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_10_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_10_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_11_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_11_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_11_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_11_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_11_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_12_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_12_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_12_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_12_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_12_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_13_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_13_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_13_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_13_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_13_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_14_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_14_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_14_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_14_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_14_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_15_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_15_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_15_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_15_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_15_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_16_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_16_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_16_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_16_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_16_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_17_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [6:0] dout_17_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_17_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire [63:0] dout_17_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_17_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  wire dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz;
  wire din_0_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_0_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_0_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_0_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_0_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_0_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_0_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_1_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_1_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_1_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_1_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_1_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_2_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_2_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_2_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_2_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_2_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_3_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_3_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_3_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_3_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_3_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_4_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_4_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_4_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_4_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_4_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_5_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_5_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_5_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_5_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_5_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_6_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_6_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_6_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_6_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_6_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_7_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_7_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_7_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_7_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_7_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_8_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_8_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_8_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_8_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_8_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_9_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_9_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_9_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_9_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_9_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_10_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_10_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_10_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_10_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_10_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_11_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_11_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_11_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_11_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_11_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_12_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_12_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_12_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_12_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_12_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_13_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_13_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_13_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_13_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_13_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_14_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_14_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_14_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_14_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_14_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_15_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_15_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_15_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_15_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_15_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_16_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_16_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_16_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_16_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_16_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_17_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [6:0] din_17_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_17_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [63:0] din_17_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_17_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire [511:0] dout_rsc_z_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  wire din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz;
  wire din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire dout_0_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_0_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_1_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_1_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_2_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_2_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_3_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_3_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_4_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_4_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_5_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_5_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_6_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_6_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_7_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_7_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_8_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_8_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_9_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_9_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_10_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_10_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_11_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_11_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_12_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_12_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_13_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_13_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_14_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_14_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_15_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_15_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_16_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_16_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud;
  wire dout_17_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud;
  wire din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud;
  wire din_17_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud;
  wire shr_mem_0_cns_R0;
  wire shr_mem_0_cns_R1;
  wire [6:0] shr_mem_0_cns_addra_shi0;
  wire [6:0] shr_mem_0_cns_addra_shi1;
  wire [6:0] shr_mem_0_cns_addrb_shi0;
  wire [6:0] shr_mem_0_cns_addrb_shi1;
  wire shr_mem_0_cns_csa_n_shi0;
  wire shr_mem_0_cns_csa_n_shi1;
  wire shr_mem_0_cns_csb_n_shi0;
  wire shr_mem_0_cns_csb_n_shi1;
  wire [63:0] shr_mem_0_cns_dinb_shi0;
  wire [63:0] shr_mem_0_cns_dinb_shi1;
  wire [63:0] shr_mem_0_cns_douta_sho0;
  wire [63:0] shr_mem_0_cns_douta_sho1;
  wire shr_mem_0_cns_unc_1;
  wire shr_mem_1_cns_R0;
  wire shr_mem_1_cns_R1;
  wire [6:0] shr_mem_1_cns_addra_shi0;
  wire [6:0] shr_mem_1_cns_addra_shi1;
  wire [6:0] shr_mem_1_cns_addrb_shi0;
  wire [6:0] shr_mem_1_cns_addrb_shi1;
  wire shr_mem_1_cns_csa_n_shi0;
  wire shr_mem_1_cns_csa_n_shi1;
  wire shr_mem_1_cns_csb_n_shi0;
  wire shr_mem_1_cns_csb_n_shi1;
  wire [63:0] shr_mem_1_cns_dinb_shi0;
  wire [63:0] shr_mem_1_cns_dinb_shi1;
  wire [63:0] shr_mem_1_cns_douta_sho0;
  wire [63:0] shr_mem_1_cns_douta_sho1;
  wire shr_mem_1_cns_unc_1;
  wire shr_mem_2_cns_R0;
  wire shr_mem_2_cns_R1;
  wire [6:0] shr_mem_2_cns_addra_shi0;
  wire [6:0] shr_mem_2_cns_addra_shi1;
  wire [6:0] shr_mem_2_cns_addrb_shi0;
  wire [6:0] shr_mem_2_cns_addrb_shi1;
  wire shr_mem_2_cns_csa_n_shi0;
  wire shr_mem_2_cns_csa_n_shi1;
  wire shr_mem_2_cns_csb_n_shi0;
  wire shr_mem_2_cns_csb_n_shi1;
  wire [63:0] shr_mem_2_cns_dinb_shi0;
  wire [63:0] shr_mem_2_cns_dinb_shi1;
  wire [63:0] shr_mem_2_cns_douta_sho0;
  wire [63:0] shr_mem_2_cns_douta_sho1;
  wire shr_mem_2_cns_unc_1;
  wire shr_mem_3_cns_R0;
  wire shr_mem_3_cns_R1;
  wire [6:0] shr_mem_3_cns_addra_shi0;
  wire [6:0] shr_mem_3_cns_addra_shi1;
  wire [6:0] shr_mem_3_cns_addrb_shi0;
  wire [6:0] shr_mem_3_cns_addrb_shi1;
  wire shr_mem_3_cns_csa_n_shi0;
  wire shr_mem_3_cns_csa_n_shi1;
  wire shr_mem_3_cns_csb_n_shi0;
  wire shr_mem_3_cns_csb_n_shi1;
  wire [63:0] shr_mem_3_cns_dinb_shi0;
  wire [63:0] shr_mem_3_cns_dinb_shi1;
  wire [63:0] shr_mem_3_cns_douta_sho0;
  wire [63:0] shr_mem_3_cns_douta_sho1;
  wire shr_mem_3_cns_unc_1;
  wire shr_mem_4_cns_R0;
  wire shr_mem_4_cns_R1;
  wire [6:0] shr_mem_4_cns_addra_shi0;
  wire [6:0] shr_mem_4_cns_addra_shi1;
  wire [6:0] shr_mem_4_cns_addrb_shi0;
  wire [6:0] shr_mem_4_cns_addrb_shi1;
  wire shr_mem_4_cns_csa_n_shi0;
  wire shr_mem_4_cns_csa_n_shi1;
  wire shr_mem_4_cns_csb_n_shi0;
  wire shr_mem_4_cns_csb_n_shi1;
  wire [63:0] shr_mem_4_cns_dinb_shi0;
  wire [63:0] shr_mem_4_cns_dinb_shi1;
  wire [63:0] shr_mem_4_cns_douta_sho0;
  wire [63:0] shr_mem_4_cns_douta_sho1;
  wire shr_mem_4_cns_unc_1;
  wire shr_mem_5_cns_R0;
  wire shr_mem_5_cns_R1;
  wire [6:0] shr_mem_5_cns_addra_shi0;
  wire [6:0] shr_mem_5_cns_addra_shi1;
  wire [6:0] shr_mem_5_cns_addrb_shi0;
  wire [6:0] shr_mem_5_cns_addrb_shi1;
  wire shr_mem_5_cns_csa_n_shi0;
  wire shr_mem_5_cns_csa_n_shi1;
  wire shr_mem_5_cns_csb_n_shi0;
  wire shr_mem_5_cns_csb_n_shi1;
  wire [63:0] shr_mem_5_cns_dinb_shi0;
  wire [63:0] shr_mem_5_cns_dinb_shi1;
  wire [63:0] shr_mem_5_cns_douta_sho0;
  wire [63:0] shr_mem_5_cns_douta_sho1;
  wire shr_mem_5_cns_unc_1;
  wire shr_mem_6_cns_R0;
  wire shr_mem_6_cns_R1;
  wire [6:0] shr_mem_6_cns_addra_shi0;
  wire [6:0] shr_mem_6_cns_addra_shi1;
  wire [6:0] shr_mem_6_cns_addrb_shi0;
  wire [6:0] shr_mem_6_cns_addrb_shi1;
  wire shr_mem_6_cns_csa_n_shi0;
  wire shr_mem_6_cns_csa_n_shi1;
  wire shr_mem_6_cns_csb_n_shi0;
  wire shr_mem_6_cns_csb_n_shi1;
  wire [63:0] shr_mem_6_cns_dinb_shi0;
  wire [63:0] shr_mem_6_cns_dinb_shi1;
  wire [63:0] shr_mem_6_cns_douta_sho0;
  wire [63:0] shr_mem_6_cns_douta_sho1;
  wire shr_mem_6_cns_unc_1;
  wire shr_mem_7_cns_R0;
  wire shr_mem_7_cns_R1;
  wire [6:0] shr_mem_7_cns_addra_shi0;
  wire [6:0] shr_mem_7_cns_addra_shi1;
  wire [6:0] shr_mem_7_cns_addrb_shi0;
  wire [6:0] shr_mem_7_cns_addrb_shi1;
  wire shr_mem_7_cns_csa_n_shi0;
  wire shr_mem_7_cns_csa_n_shi1;
  wire shr_mem_7_cns_csb_n_shi0;
  wire shr_mem_7_cns_csb_n_shi1;
  wire [63:0] shr_mem_7_cns_dinb_shi0;
  wire [63:0] shr_mem_7_cns_dinb_shi1;
  wire [63:0] shr_mem_7_cns_douta_sho0;
  wire [63:0] shr_mem_7_cns_douta_sho1;
  wire shr_mem_7_cns_unc_1;
  wire shr_mem_8_cns_R0;
  wire shr_mem_8_cns_R1;
  wire [6:0] shr_mem_8_cns_addra_shi0;
  wire [6:0] shr_mem_8_cns_addra_shi1;
  wire [6:0] shr_mem_8_cns_addrb_shi0;
  wire [6:0] shr_mem_8_cns_addrb_shi1;
  wire shr_mem_8_cns_csa_n_shi0;
  wire shr_mem_8_cns_csa_n_shi1;
  wire shr_mem_8_cns_csb_n_shi0;
  wire shr_mem_8_cns_csb_n_shi1;
  wire [63:0] shr_mem_8_cns_dinb_shi0;
  wire [63:0] shr_mem_8_cns_dinb_shi1;
  wire [63:0] shr_mem_8_cns_douta_sho0;
  wire [63:0] shr_mem_8_cns_douta_sho1;
  wire shr_mem_8_cns_unc_1;
  wire shr_mem_9_cns_R0;
  wire shr_mem_9_cns_R1;
  wire [6:0] shr_mem_9_cns_addra_shi0;
  wire [6:0] shr_mem_9_cns_addra_shi1;
  wire [6:0] shr_mem_9_cns_addrb_shi0;
  wire [6:0] shr_mem_9_cns_addrb_shi1;
  wire shr_mem_9_cns_csa_n_shi0;
  wire shr_mem_9_cns_csa_n_shi1;
  wire shr_mem_9_cns_csb_n_shi0;
  wire shr_mem_9_cns_csb_n_shi1;
  wire [63:0] shr_mem_9_cns_dinb_shi0;
  wire [63:0] shr_mem_9_cns_dinb_shi1;
  wire [63:0] shr_mem_9_cns_douta_sho0;
  wire [63:0] shr_mem_9_cns_douta_sho1;
  wire shr_mem_9_cns_unc_1;
  wire shr_mem_10_cns_R0;
  wire shr_mem_10_cns_R1;
  wire [6:0] shr_mem_10_cns_addra_shi0;
  wire [6:0] shr_mem_10_cns_addra_shi1;
  wire [6:0] shr_mem_10_cns_addrb_shi0;
  wire [6:0] shr_mem_10_cns_addrb_shi1;
  wire shr_mem_10_cns_csa_n_shi0;
  wire shr_mem_10_cns_csa_n_shi1;
  wire shr_mem_10_cns_csb_n_shi0;
  wire shr_mem_10_cns_csb_n_shi1;
  wire [63:0] shr_mem_10_cns_dinb_shi0;
  wire [63:0] shr_mem_10_cns_dinb_shi1;
  wire [63:0] shr_mem_10_cns_douta_sho0;
  wire [63:0] shr_mem_10_cns_douta_sho1;
  wire shr_mem_10_cns_unc_1;
  wire shr_mem_11_cns_R0;
  wire shr_mem_11_cns_R1;
  wire [6:0] shr_mem_11_cns_addra_shi0;
  wire [6:0] shr_mem_11_cns_addra_shi1;
  wire [6:0] shr_mem_11_cns_addrb_shi0;
  wire [6:0] shr_mem_11_cns_addrb_shi1;
  wire shr_mem_11_cns_csa_n_shi0;
  wire shr_mem_11_cns_csa_n_shi1;
  wire shr_mem_11_cns_csb_n_shi0;
  wire shr_mem_11_cns_csb_n_shi1;
  wire [63:0] shr_mem_11_cns_dinb_shi0;
  wire [63:0] shr_mem_11_cns_dinb_shi1;
  wire [63:0] shr_mem_11_cns_douta_sho0;
  wire [63:0] shr_mem_11_cns_douta_sho1;
  wire shr_mem_11_cns_unc_1;
  wire shr_mem_12_cns_R0;
  wire shr_mem_12_cns_R1;
  wire [6:0] shr_mem_12_cns_addra_shi0;
  wire [6:0] shr_mem_12_cns_addra_shi1;
  wire [6:0] shr_mem_12_cns_addrb_shi0;
  wire [6:0] shr_mem_12_cns_addrb_shi1;
  wire shr_mem_12_cns_csa_n_shi0;
  wire shr_mem_12_cns_csa_n_shi1;
  wire shr_mem_12_cns_csb_n_shi0;
  wire shr_mem_12_cns_csb_n_shi1;
  wire [63:0] shr_mem_12_cns_dinb_shi0;
  wire [63:0] shr_mem_12_cns_dinb_shi1;
  wire [63:0] shr_mem_12_cns_douta_sho0;
  wire [63:0] shr_mem_12_cns_douta_sho1;
  wire shr_mem_12_cns_unc_1;
  wire shr_mem_13_cns_R0;
  wire shr_mem_13_cns_R1;
  wire [6:0] shr_mem_13_cns_addra_shi0;
  wire [6:0] shr_mem_13_cns_addra_shi1;
  wire [6:0] shr_mem_13_cns_addrb_shi0;
  wire [6:0] shr_mem_13_cns_addrb_shi1;
  wire shr_mem_13_cns_csa_n_shi0;
  wire shr_mem_13_cns_csa_n_shi1;
  wire shr_mem_13_cns_csb_n_shi0;
  wire shr_mem_13_cns_csb_n_shi1;
  wire [63:0] shr_mem_13_cns_dinb_shi0;
  wire [63:0] shr_mem_13_cns_dinb_shi1;
  wire [63:0] shr_mem_13_cns_douta_sho0;
  wire [63:0] shr_mem_13_cns_douta_sho1;
  wire shr_mem_13_cns_unc_1;
  wire shr_mem_14_cns_R0;
  wire shr_mem_14_cns_R1;
  wire [6:0] shr_mem_14_cns_addra_shi0;
  wire [6:0] shr_mem_14_cns_addra_shi1;
  wire [6:0] shr_mem_14_cns_addrb_shi0;
  wire [6:0] shr_mem_14_cns_addrb_shi1;
  wire shr_mem_14_cns_csa_n_shi0;
  wire shr_mem_14_cns_csa_n_shi1;
  wire shr_mem_14_cns_csb_n_shi0;
  wire shr_mem_14_cns_csb_n_shi1;
  wire [63:0] shr_mem_14_cns_dinb_shi0;
  wire [63:0] shr_mem_14_cns_dinb_shi1;
  wire [63:0] shr_mem_14_cns_douta_sho0;
  wire [63:0] shr_mem_14_cns_douta_sho1;
  wire shr_mem_14_cns_unc_1;
  wire shr_mem_15_cns_R0;
  wire shr_mem_15_cns_R1;
  wire [6:0] shr_mem_15_cns_addra_shi0;
  wire [6:0] shr_mem_15_cns_addra_shi1;
  wire [6:0] shr_mem_15_cns_addrb_shi0;
  wire [6:0] shr_mem_15_cns_addrb_shi1;
  wire shr_mem_15_cns_csa_n_shi0;
  wire shr_mem_15_cns_csa_n_shi1;
  wire shr_mem_15_cns_csb_n_shi0;
  wire shr_mem_15_cns_csb_n_shi1;
  wire [63:0] shr_mem_15_cns_dinb_shi0;
  wire [63:0] shr_mem_15_cns_dinb_shi1;
  wire [63:0] shr_mem_15_cns_douta_sho0;
  wire [63:0] shr_mem_15_cns_douta_sho1;
  wire shr_mem_15_cns_unc_1;
  wire shr_mem_16_cns_R0;
  wire shr_mem_16_cns_R1;
  wire [6:0] shr_mem_16_cns_addra_shi0;
  wire [6:0] shr_mem_16_cns_addra_shi1;
  wire [6:0] shr_mem_16_cns_addrb_shi0;
  wire [6:0] shr_mem_16_cns_addrb_shi1;
  wire shr_mem_16_cns_csa_n_shi0;
  wire shr_mem_16_cns_csa_n_shi1;
  wire shr_mem_16_cns_csb_n_shi0;
  wire shr_mem_16_cns_csb_n_shi1;
  wire [63:0] shr_mem_16_cns_dinb_shi0;
  wire [63:0] shr_mem_16_cns_dinb_shi1;
  wire [63:0] shr_mem_16_cns_douta_sho0;
  wire [63:0] shr_mem_16_cns_douta_sho1;
  wire shr_mem_16_cns_unc_1;
  wire shr_mem_17_cns_R0;
  wire shr_mem_17_cns_R1;
  wire [6:0] shr_mem_17_cns_addra_shi0;
  wire [6:0] shr_mem_17_cns_addra_shi1;
  wire [6:0] shr_mem_17_cns_addrb_shi0;
  wire [6:0] shr_mem_17_cns_addrb_shi1;
  wire shr_mem_17_cns_csa_n_shi0;
  wire shr_mem_17_cns_csa_n_shi1;
  wire shr_mem_17_cns_csb_n_shi0;
  wire shr_mem_17_cns_csb_n_shi1;
  wire [63:0] shr_mem_17_cns_dinb_shi0;
  wire [63:0] shr_mem_17_cns_dinb_shi1;
  wire [63:0] shr_mem_17_cns_douta_sho0;
  wire [63:0] shr_mem_17_cns_douta_sho1;
  wire shr_mem_17_cns_unc_1;
  wire shr_mem_0_cns_S1_iff;
  wire shr_mem_0_cns_S0_iff;
  wire shr_mem_1_cns_S1_iff;
  wire din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_1_cns_S0_iff;
  wire shr_mem_2_cns_S1_iff;
  wire din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_2_cns_S0_iff;
  wire shr_mem_3_cns_S1_iff;
  wire din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_3_cns_S0_iff;
  wire shr_mem_4_cns_S1_iff;
  wire din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_4_cns_S0_iff;
  wire shr_mem_5_cns_S1_iff;
  wire din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_5_cns_S0_iff;
  wire shr_mem_6_cns_S1_iff;
  wire din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_6_cns_S0_iff;
  wire shr_mem_7_cns_S1_iff;
  wire din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_7_cns_S0_iff;
  wire shr_mem_8_cns_S1_iff;
  wire din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_8_cns_S0_iff;
  wire shr_mem_9_cns_S1_iff;
  wire din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_9_cns_S0_iff;
  wire shr_mem_10_cns_S1_iff;
  wire din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_10_cns_S0_iff;
  wire shr_mem_11_cns_S1_iff;
  wire din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_11_cns_S0_iff;
  wire shr_mem_12_cns_S1_iff;
  wire din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_12_cns_S0_iff;
  wire shr_mem_13_cns_S1_iff;
  wire din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_13_cns_S0_iff;
  wire shr_mem_14_cns_S1_iff;
  wire din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_14_cns_S0_iff;
  wire shr_mem_15_cns_S1_iff;
  wire din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_15_cns_S0_iff;
  wire shr_mem_16_cns_S1_iff;
  wire din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_16_cns_S0_iff;
  wire shr_mem_17_cns_S1_iff;
  wire din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff;
  wire din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff;
  wire dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff;
  wire dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff;
  wire shr_mem_17_cns_S0_iff;
  wire shr_mem_0_cns_S0_dmo;
  wire shr_mem_0_cns_S1_dmo;
  wire shr_mem_1_cns_S0_dmo;
  wire shr_mem_1_cns_S1_dmo;
  wire shr_mem_2_cns_S0_dmo;
  wire shr_mem_2_cns_S1_dmo;
  wire shr_mem_3_cns_S0_dmo;
  wire shr_mem_3_cns_S1_dmo;
  wire shr_mem_4_cns_S0_dmo;
  wire shr_mem_4_cns_S1_dmo;
  wire shr_mem_5_cns_S0_dmo;
  wire shr_mem_5_cns_S1_dmo;
  wire shr_mem_6_cns_S0_dmo;
  wire shr_mem_6_cns_S1_dmo;
  wire shr_mem_7_cns_S0_dmo;
  wire shr_mem_7_cns_S1_dmo;
  wire shr_mem_8_cns_S0_dmo;
  wire shr_mem_8_cns_S1_dmo;
  wire shr_mem_9_cns_S0_dmo;
  wire shr_mem_9_cns_S1_dmo;
  wire shr_mem_10_cns_S0_dmo;
  wire shr_mem_10_cns_S1_dmo;
  wire shr_mem_11_cns_S0_dmo;
  wire shr_mem_11_cns_S1_dmo;
  wire shr_mem_12_cns_S0_dmo;
  wire shr_mem_12_cns_S1_dmo;
  wire shr_mem_13_cns_S0_dmo;
  wire shr_mem_13_cns_S1_dmo;
  wire shr_mem_14_cns_S0_dmo;
  wire shr_mem_14_cns_S1_dmo;
  wire shr_mem_15_cns_S0_dmo;
  wire shr_mem_15_cns_S1_dmo;
  wire shr_mem_16_cns_S0_dmo;
  wire shr_mem_16_cns_S1_dmo;
  wire shr_mem_17_cns_S0_dmo;
  wire shr_mem_17_cns_S1_dmo;


  // Interconnect Declarations for Component Instantiations 
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_0_cns_comp (
      .addra(shr_mem_0_cns_addra_shi0),
      .addrb(shr_mem_0_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_0_cns_csa_n_shi0),
      .csb_n(shr_mem_0_cns_csb_n_shi0),
      .dinb(shr_mem_0_cns_dinb_shi0),
      .douta(shr_mem_0_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_0_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_0_cns_comp_1 (
      .addra(shr_mem_0_cns_addra_shi1),
      .addrb(shr_mem_0_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_0_cns_csa_n_shi1),
      .csb_n(shr_mem_0_cns_csb_n_shi1),
      .dinb(shr_mem_0_cns_dinb_shi1),
      .douta(shr_mem_0_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_0_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_1_cns_comp (
      .addra(shr_mem_1_cns_addra_shi0),
      .addrb(shr_mem_1_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_1_cns_csa_n_shi0),
      .csb_n(shr_mem_1_cns_csb_n_shi0),
      .dinb(shr_mem_1_cns_dinb_shi0),
      .douta(shr_mem_1_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_1_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_1_cns_comp_1 (
      .addra(shr_mem_1_cns_addra_shi1),
      .addrb(shr_mem_1_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_1_cns_csa_n_shi1),
      .csb_n(shr_mem_1_cns_csb_n_shi1),
      .dinb(shr_mem_1_cns_dinb_shi1),
      .douta(shr_mem_1_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_1_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_2_cns_comp (
      .addra(shr_mem_2_cns_addra_shi0),
      .addrb(shr_mem_2_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_2_cns_csa_n_shi0),
      .csb_n(shr_mem_2_cns_csb_n_shi0),
      .dinb(shr_mem_2_cns_dinb_shi0),
      .douta(shr_mem_2_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_2_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_2_cns_comp_1 (
      .addra(shr_mem_2_cns_addra_shi1),
      .addrb(shr_mem_2_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_2_cns_csa_n_shi1),
      .csb_n(shr_mem_2_cns_csb_n_shi1),
      .dinb(shr_mem_2_cns_dinb_shi1),
      .douta(shr_mem_2_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_2_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_3_cns_comp (
      .addra(shr_mem_3_cns_addra_shi0),
      .addrb(shr_mem_3_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_3_cns_csa_n_shi0),
      .csb_n(shr_mem_3_cns_csb_n_shi0),
      .dinb(shr_mem_3_cns_dinb_shi0),
      .douta(shr_mem_3_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_3_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_3_cns_comp_1 (
      .addra(shr_mem_3_cns_addra_shi1),
      .addrb(shr_mem_3_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_3_cns_csa_n_shi1),
      .csb_n(shr_mem_3_cns_csb_n_shi1),
      .dinb(shr_mem_3_cns_dinb_shi1),
      .douta(shr_mem_3_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_3_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_4_cns_comp (
      .addra(shr_mem_4_cns_addra_shi0),
      .addrb(shr_mem_4_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_4_cns_csa_n_shi0),
      .csb_n(shr_mem_4_cns_csb_n_shi0),
      .dinb(shr_mem_4_cns_dinb_shi0),
      .douta(shr_mem_4_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_4_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_4_cns_comp_1 (
      .addra(shr_mem_4_cns_addra_shi1),
      .addrb(shr_mem_4_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_4_cns_csa_n_shi1),
      .csb_n(shr_mem_4_cns_csb_n_shi1),
      .dinb(shr_mem_4_cns_dinb_shi1),
      .douta(shr_mem_4_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_4_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_5_cns_comp (
      .addra(shr_mem_5_cns_addra_shi0),
      .addrb(shr_mem_5_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_5_cns_csa_n_shi0),
      .csb_n(shr_mem_5_cns_csb_n_shi0),
      .dinb(shr_mem_5_cns_dinb_shi0),
      .douta(shr_mem_5_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_5_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_5_cns_comp_1 (
      .addra(shr_mem_5_cns_addra_shi1),
      .addrb(shr_mem_5_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_5_cns_csa_n_shi1),
      .csb_n(shr_mem_5_cns_csb_n_shi1),
      .dinb(shr_mem_5_cns_dinb_shi1),
      .douta(shr_mem_5_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_5_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_6_cns_comp (
      .addra(shr_mem_6_cns_addra_shi0),
      .addrb(shr_mem_6_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_6_cns_csa_n_shi0),
      .csb_n(shr_mem_6_cns_csb_n_shi0),
      .dinb(shr_mem_6_cns_dinb_shi0),
      .douta(shr_mem_6_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_6_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_6_cns_comp_1 (
      .addra(shr_mem_6_cns_addra_shi1),
      .addrb(shr_mem_6_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_6_cns_csa_n_shi1),
      .csb_n(shr_mem_6_cns_csb_n_shi1),
      .dinb(shr_mem_6_cns_dinb_shi1),
      .douta(shr_mem_6_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_6_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_7_cns_comp (
      .addra(shr_mem_7_cns_addra_shi0),
      .addrb(shr_mem_7_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_7_cns_csa_n_shi0),
      .csb_n(shr_mem_7_cns_csb_n_shi0),
      .dinb(shr_mem_7_cns_dinb_shi0),
      .douta(shr_mem_7_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_7_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_7_cns_comp_1 (
      .addra(shr_mem_7_cns_addra_shi1),
      .addrb(shr_mem_7_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_7_cns_csa_n_shi1),
      .csb_n(shr_mem_7_cns_csb_n_shi1),
      .dinb(shr_mem_7_cns_dinb_shi1),
      .douta(shr_mem_7_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_7_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_8_cns_comp (
      .addra(shr_mem_8_cns_addra_shi0),
      .addrb(shr_mem_8_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_8_cns_csa_n_shi0),
      .csb_n(shr_mem_8_cns_csb_n_shi0),
      .dinb(shr_mem_8_cns_dinb_shi0),
      .douta(shr_mem_8_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_8_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_8_cns_comp_1 (
      .addra(shr_mem_8_cns_addra_shi1),
      .addrb(shr_mem_8_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_8_cns_csa_n_shi1),
      .csb_n(shr_mem_8_cns_csb_n_shi1),
      .dinb(shr_mem_8_cns_dinb_shi1),
      .douta(shr_mem_8_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_8_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_9_cns_comp (
      .addra(shr_mem_9_cns_addra_shi0),
      .addrb(shr_mem_9_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_9_cns_csa_n_shi0),
      .csb_n(shr_mem_9_cns_csb_n_shi0),
      .dinb(shr_mem_9_cns_dinb_shi0),
      .douta(shr_mem_9_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_9_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_9_cns_comp_1 (
      .addra(shr_mem_9_cns_addra_shi1),
      .addrb(shr_mem_9_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_9_cns_csa_n_shi1),
      .csb_n(shr_mem_9_cns_csb_n_shi1),
      .dinb(shr_mem_9_cns_dinb_shi1),
      .douta(shr_mem_9_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_9_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_10_cns_comp (
      .addra(shr_mem_10_cns_addra_shi0),
      .addrb(shr_mem_10_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_10_cns_csa_n_shi0),
      .csb_n(shr_mem_10_cns_csb_n_shi0),
      .dinb(shr_mem_10_cns_dinb_shi0),
      .douta(shr_mem_10_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_10_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_10_cns_comp_1 (
      .addra(shr_mem_10_cns_addra_shi1),
      .addrb(shr_mem_10_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_10_cns_csa_n_shi1),
      .csb_n(shr_mem_10_cns_csb_n_shi1),
      .dinb(shr_mem_10_cns_dinb_shi1),
      .douta(shr_mem_10_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_10_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_11_cns_comp (
      .addra(shr_mem_11_cns_addra_shi0),
      .addrb(shr_mem_11_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_11_cns_csa_n_shi0),
      .csb_n(shr_mem_11_cns_csb_n_shi0),
      .dinb(shr_mem_11_cns_dinb_shi0),
      .douta(shr_mem_11_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_11_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_11_cns_comp_1 (
      .addra(shr_mem_11_cns_addra_shi1),
      .addrb(shr_mem_11_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_11_cns_csa_n_shi1),
      .csb_n(shr_mem_11_cns_csb_n_shi1),
      .dinb(shr_mem_11_cns_dinb_shi1),
      .douta(shr_mem_11_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_11_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_12_cns_comp (
      .addra(shr_mem_12_cns_addra_shi0),
      .addrb(shr_mem_12_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_12_cns_csa_n_shi0),
      .csb_n(shr_mem_12_cns_csb_n_shi0),
      .dinb(shr_mem_12_cns_dinb_shi0),
      .douta(shr_mem_12_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_12_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_12_cns_comp_1 (
      .addra(shr_mem_12_cns_addra_shi1),
      .addrb(shr_mem_12_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_12_cns_csa_n_shi1),
      .csb_n(shr_mem_12_cns_csb_n_shi1),
      .dinb(shr_mem_12_cns_dinb_shi1),
      .douta(shr_mem_12_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_12_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_13_cns_comp (
      .addra(shr_mem_13_cns_addra_shi0),
      .addrb(shr_mem_13_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_13_cns_csa_n_shi0),
      .csb_n(shr_mem_13_cns_csb_n_shi0),
      .dinb(shr_mem_13_cns_dinb_shi0),
      .douta(shr_mem_13_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_13_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_13_cns_comp_1 (
      .addra(shr_mem_13_cns_addra_shi1),
      .addrb(shr_mem_13_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_13_cns_csa_n_shi1),
      .csb_n(shr_mem_13_cns_csb_n_shi1),
      .dinb(shr_mem_13_cns_dinb_shi1),
      .douta(shr_mem_13_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_13_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_14_cns_comp (
      .addra(shr_mem_14_cns_addra_shi0),
      .addrb(shr_mem_14_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_14_cns_csa_n_shi0),
      .csb_n(shr_mem_14_cns_csb_n_shi0),
      .dinb(shr_mem_14_cns_dinb_shi0),
      .douta(shr_mem_14_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_14_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_14_cns_comp_1 (
      .addra(shr_mem_14_cns_addra_shi1),
      .addrb(shr_mem_14_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_14_cns_csa_n_shi1),
      .csb_n(shr_mem_14_cns_csb_n_shi1),
      .dinb(shr_mem_14_cns_dinb_shi1),
      .douta(shr_mem_14_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_14_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_15_cns_comp (
      .addra(shr_mem_15_cns_addra_shi0),
      .addrb(shr_mem_15_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_15_cns_csa_n_shi0),
      .csb_n(shr_mem_15_cns_csb_n_shi0),
      .dinb(shr_mem_15_cns_dinb_shi0),
      .douta(shr_mem_15_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_15_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_15_cns_comp_1 (
      .addra(shr_mem_15_cns_addra_shi1),
      .addrb(shr_mem_15_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_15_cns_csa_n_shi1),
      .csb_n(shr_mem_15_cns_csb_n_shi1),
      .dinb(shr_mem_15_cns_dinb_shi1),
      .douta(shr_mem_15_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_15_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_16_cns_comp (
      .addra(shr_mem_16_cns_addra_shi0),
      .addrb(shr_mem_16_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_16_cns_csa_n_shi0),
      .csb_n(shr_mem_16_cns_csb_n_shi0),
      .dinb(shr_mem_16_cns_dinb_shi0),
      .douta(shr_mem_16_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_16_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_16_cns_comp_1 (
      .addra(shr_mem_16_cns_addra_shi1),
      .addrb(shr_mem_16_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_16_cns_csa_n_shi1),
      .csb_n(shr_mem_16_cns_csb_n_shi1),
      .dinb(shr_mem_16_cns_dinb_shi1),
      .douta(shr_mem_16_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_16_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_17_cns_comp (
      .addra(shr_mem_17_cns_addra_shi0),
      .addrb(shr_mem_17_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_17_cns_csa_n_shi0),
      .csb_n(shr_mem_17_cns_csb_n_shi0),
      .dinb(shr_mem_17_cns_dinb_shi0),
      .douta(shr_mem_17_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_17_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_17_cns_comp_1 (
      .addra(shr_mem_17_cns_addra_shi1),
      .addrb(shr_mem_17_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_17_cns_csa_n_shi1),
      .csb_n(shr_mem_17_cns_csb_n_shi1),
      .dinb(shr_mem_17_cns_dinb_shi1),
      .douta(shr_mem_17_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_17_cns_unc_1)
    );
  WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_1 WRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(din_rsc_z),
      .din_rsc_vz(din_rsc_vz),
      .din_rsc_lz(din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_0_rsc_csa_n(dout_0_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_csb_n(dout_0_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_addra(dout_0_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_addrb(dout_0_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_dinb(dout_0_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_douta(dout_0_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_req_vz(dout_0_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_rls_lz(dout_0_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_1_rsc_csa_n(dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_csb_n(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_addra(dout_1_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_addrb(dout_1_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_dinb(dout_1_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_douta(dout_1_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_req_vz(dout_1_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_rls_lz(dout_1_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_2_rsc_csa_n(dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_csb_n(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_addra(dout_2_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_addrb(dout_2_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_dinb(dout_2_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_douta(dout_2_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_req_vz(dout_2_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_rls_lz(dout_2_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_3_rsc_csa_n(dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_csb_n(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_addra(dout_3_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_addrb(dout_3_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_dinb(dout_3_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_douta(dout_3_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_req_vz(dout_3_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_rls_lz(dout_3_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_4_rsc_csa_n(dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_csb_n(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_addra(dout_4_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_addrb(dout_4_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_dinb(dout_4_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_douta(dout_4_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_req_vz(dout_4_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_rls_lz(dout_4_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_5_rsc_csa_n(dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_csb_n(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_addra(dout_5_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_addrb(dout_5_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_dinb(dout_5_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_douta(dout_5_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_req_vz(dout_5_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_rls_lz(dout_5_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_6_rsc_csa_n(dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_csb_n(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_addra(dout_6_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_addrb(dout_6_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_dinb(dout_6_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_douta(dout_6_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_req_vz(dout_6_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_rls_lz(dout_6_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_7_rsc_csa_n(dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_csb_n(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_addra(dout_7_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_addrb(dout_7_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_dinb(dout_7_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_douta(dout_7_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_req_vz(dout_7_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_rls_lz(dout_7_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_8_rsc_csa_n(dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_csb_n(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_addra(dout_8_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_addrb(dout_8_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_dinb(dout_8_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_douta(dout_8_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_req_vz(dout_8_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_rls_lz(dout_8_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_9_rsc_csa_n(dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_csb_n(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_addra(dout_9_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_addrb(dout_9_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_dinb(dout_9_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_douta(dout_9_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_req_vz(dout_9_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_rls_lz(dout_9_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_10_rsc_csa_n(dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_csb_n(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_addra(dout_10_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_addrb(dout_10_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_dinb(dout_10_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_douta(dout_10_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_req_vz(dout_10_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_rls_lz(dout_10_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_11_rsc_csa_n(dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_csb_n(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_addra(dout_11_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_addrb(dout_11_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_dinb(dout_11_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_douta(dout_11_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_req_vz(dout_11_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_rls_lz(dout_11_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_12_rsc_csa_n(dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_csb_n(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_addra(dout_12_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_addrb(dout_12_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_dinb(dout_12_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_douta(dout_12_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_req_vz(dout_12_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_rls_lz(dout_12_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_13_rsc_csa_n(dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_csb_n(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_addra(dout_13_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_addrb(dout_13_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_dinb(dout_13_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_douta(dout_13_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_req_vz(dout_13_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_rls_lz(dout_13_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_14_rsc_csa_n(dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_csb_n(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_addra(dout_14_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_addrb(dout_14_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_dinb(dout_14_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_douta(dout_14_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_req_vz(dout_14_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_rls_lz(dout_14_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_15_rsc_csa_n(dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_csb_n(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_addra(dout_15_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_addrb(dout_15_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_dinb(dout_15_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_douta(dout_15_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_req_vz(dout_15_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_rls_lz(dout_15_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_16_rsc_csa_n(dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_csb_n(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_addra(dout_16_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_addrb(dout_16_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_dinb(dout_16_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_douta(dout_16_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_req_vz(dout_16_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_rls_lz(dout_16_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_17_rsc_csa_n(dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_csb_n(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_addra(dout_17_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_addrb(dout_17_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_dinb(dout_17_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_douta(dout_17_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_req_vz(dout_17_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_rls_lz(dout_17_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .clamp_mem(clamp_mem),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n)
    );
  READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_1 READ_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst (
      .clk(clk),
      .rst(rst),
      .din_0_rsc_csa_n(din_0_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_csb_n(din_0_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_addra(din_0_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_addrb(din_0_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_dinb(din_0_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_douta(din_0_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_req_vz(din_0_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_rls_lz(din_0_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_1_rsc_csa_n(din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_csb_n(din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_addra(din_1_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_addrb(din_1_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_dinb(din_1_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_douta(din_1_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_req_vz(din_1_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_rls_lz(din_1_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_2_rsc_csa_n(din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_csb_n(din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_addra(din_2_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_addrb(din_2_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_dinb(din_2_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_douta(din_2_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_req_vz(din_2_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_rls_lz(din_2_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_3_rsc_csa_n(din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_csb_n(din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_addra(din_3_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_addrb(din_3_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_dinb(din_3_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_douta(din_3_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_req_vz(din_3_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_rls_lz(din_3_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_4_rsc_csa_n(din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_csb_n(din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_addra(din_4_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_addrb(din_4_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_dinb(din_4_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_douta(din_4_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_req_vz(din_4_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_rls_lz(din_4_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_5_rsc_csa_n(din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_csb_n(din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_addra(din_5_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_addrb(din_5_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_dinb(din_5_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_douta(din_5_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_req_vz(din_5_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_rls_lz(din_5_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_6_rsc_csa_n(din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_csb_n(din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_addra(din_6_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_addrb(din_6_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_dinb(din_6_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_douta(din_6_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_req_vz(din_6_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_rls_lz(din_6_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_7_rsc_csa_n(din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_csb_n(din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_addra(din_7_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_addrb(din_7_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_dinb(din_7_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_douta(din_7_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_req_vz(din_7_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_rls_lz(din_7_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_8_rsc_csa_n(din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_csb_n(din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_addra(din_8_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_addrb(din_8_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_dinb(din_8_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_douta(din_8_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_req_vz(din_8_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_rls_lz(din_8_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_9_rsc_csa_n(din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_csb_n(din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_addra(din_9_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_addrb(din_9_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_dinb(din_9_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_douta(din_9_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_req_vz(din_9_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_rls_lz(din_9_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_10_rsc_csa_n(din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_csb_n(din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_addra(din_10_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_addrb(din_10_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_dinb(din_10_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_douta(din_10_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_req_vz(din_10_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_rls_lz(din_10_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_11_rsc_csa_n(din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_csb_n(din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_addra(din_11_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_addrb(din_11_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_dinb(din_11_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_douta(din_11_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_req_vz(din_11_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_rls_lz(din_11_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_12_rsc_csa_n(din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_csb_n(din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_addra(din_12_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_addrb(din_12_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_dinb(din_12_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_douta(din_12_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_req_vz(din_12_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_rls_lz(din_12_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_13_rsc_csa_n(din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_csb_n(din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_addra(din_13_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_addrb(din_13_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_dinb(din_13_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_douta(din_13_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_req_vz(din_13_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_rls_lz(din_13_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_14_rsc_csa_n(din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_csb_n(din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_addra(din_14_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_addrb(din_14_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_dinb(din_14_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_douta(din_14_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_req_vz(din_14_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_rls_lz(din_14_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_15_rsc_csa_n(din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_csb_n(din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_addra(din_15_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_addrb(din_15_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_dinb(din_15_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_douta(din_15_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_req_vz(din_15_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_rls_lz(din_15_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_16_rsc_csa_n(din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_csb_n(din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_addra(din_16_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_addrb(din_16_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_dinb(din_16_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_douta(din_16_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_req_vz(din_16_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_rls_lz(din_16_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .din_17_rsc_csa_n(din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_csb_n(din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_addra(din_17_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_addrb(din_17_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_dinb(din_17_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_douta(din_17_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_req_vz(din_17_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_rls_lz(din_17_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .dout_rsc_z(dout_rsc_z_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .dout_rsc_vz(dout_rsc_vz),
      .dout_rsc_lz(dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud)
    );
  unreg_hier_69 unreg (
      .in_0(shr_mem_0_cns_S0_iff),
      .out_0(shr_mem_0_cns_R0)
    );
  unreg_hier_69 unreg_1 (
      .in_0(shr_mem_0_cns_S1_iff),
      .out_0(shr_mem_0_cns_R1)
    );
  unreg_hier_69 unreg_2 (
      .in_0(shr_mem_1_cns_S0_iff),
      .out_0(shr_mem_1_cns_R0)
    );
  unreg_hier_69 unreg_3 (
      .in_0(shr_mem_1_cns_S1_iff),
      .out_0(shr_mem_1_cns_R1)
    );
  unreg_hier_69 unreg_4 (
      .in_0(shr_mem_2_cns_S0_iff),
      .out_0(shr_mem_2_cns_R0)
    );
  unreg_hier_69 unreg_5 (
      .in_0(shr_mem_2_cns_S1_iff),
      .out_0(shr_mem_2_cns_R1)
    );
  unreg_hier_69 unreg_6 (
      .in_0(shr_mem_3_cns_S0_iff),
      .out_0(shr_mem_3_cns_R0)
    );
  unreg_hier_69 unreg_7 (
      .in_0(shr_mem_3_cns_S1_iff),
      .out_0(shr_mem_3_cns_R1)
    );
  unreg_hier_69 unreg_8 (
      .in_0(shr_mem_4_cns_S0_iff),
      .out_0(shr_mem_4_cns_R0)
    );
  unreg_hier_69 unreg_9 (
      .in_0(shr_mem_4_cns_S1_iff),
      .out_0(shr_mem_4_cns_R1)
    );
  unreg_hier_69 unreg_10 (
      .in_0(shr_mem_5_cns_S0_iff),
      .out_0(shr_mem_5_cns_R0)
    );
  unreg_hier_69 unreg_11 (
      .in_0(shr_mem_5_cns_S1_iff),
      .out_0(shr_mem_5_cns_R1)
    );
  unreg_hier_69 unreg_12 (
      .in_0(shr_mem_6_cns_S0_iff),
      .out_0(shr_mem_6_cns_R0)
    );
  unreg_hier_69 unreg_13 (
      .in_0(shr_mem_6_cns_S1_iff),
      .out_0(shr_mem_6_cns_R1)
    );
  unreg_hier_69 unreg_14 (
      .in_0(shr_mem_7_cns_S0_iff),
      .out_0(shr_mem_7_cns_R0)
    );
  unreg_hier_69 unreg_15 (
      .in_0(shr_mem_7_cns_S1_iff),
      .out_0(shr_mem_7_cns_R1)
    );
  unreg_hier_69 unreg_16 (
      .in_0(shr_mem_8_cns_S0_iff),
      .out_0(shr_mem_8_cns_R0)
    );
  unreg_hier_69 unreg_17 (
      .in_0(shr_mem_8_cns_S1_iff),
      .out_0(shr_mem_8_cns_R1)
    );
  unreg_hier_69 unreg_18 (
      .in_0(shr_mem_9_cns_S0_iff),
      .out_0(shr_mem_9_cns_R0)
    );
  unreg_hier_69 unreg_19 (
      .in_0(shr_mem_9_cns_S1_iff),
      .out_0(shr_mem_9_cns_R1)
    );
  unreg_hier_69 unreg_20 (
      .in_0(shr_mem_10_cns_S0_iff),
      .out_0(shr_mem_10_cns_R0)
    );
  unreg_hier_69 unreg_21 (
      .in_0(shr_mem_10_cns_S1_iff),
      .out_0(shr_mem_10_cns_R1)
    );
  unreg_hier_69 unreg_22 (
      .in_0(shr_mem_11_cns_S0_iff),
      .out_0(shr_mem_11_cns_R0)
    );
  unreg_hier_69 unreg_23 (
      .in_0(shr_mem_11_cns_S1_iff),
      .out_0(shr_mem_11_cns_R1)
    );
  unreg_hier_69 unreg_24 (
      .in_0(shr_mem_12_cns_S0_iff),
      .out_0(shr_mem_12_cns_R0)
    );
  unreg_hier_69 unreg_25 (
      .in_0(shr_mem_12_cns_S1_iff),
      .out_0(shr_mem_12_cns_R1)
    );
  unreg_hier_69 unreg_26 (
      .in_0(shr_mem_13_cns_S0_iff),
      .out_0(shr_mem_13_cns_R0)
    );
  unreg_hier_69 unreg_27 (
      .in_0(shr_mem_13_cns_S1_iff),
      .out_0(shr_mem_13_cns_R1)
    );
  unreg_hier_69 unreg_28 (
      .in_0(shr_mem_14_cns_S0_iff),
      .out_0(shr_mem_14_cns_R0)
    );
  unreg_hier_69 unreg_29 (
      .in_0(shr_mem_14_cns_S1_iff),
      .out_0(shr_mem_14_cns_R1)
    );
  unreg_hier_69 unreg_30 (
      .in_0(shr_mem_15_cns_S0_iff),
      .out_0(shr_mem_15_cns_R0)
    );
  unreg_hier_69 unreg_31 (
      .in_0(shr_mem_15_cns_S1_iff),
      .out_0(shr_mem_15_cns_R1)
    );
  unreg_hier_69 unreg_32 (
      .in_0(shr_mem_16_cns_S0_iff),
      .out_0(shr_mem_16_cns_R0)
    );
  unreg_hier_69 unreg_33 (
      .in_0(shr_mem_16_cns_S1_iff),
      .out_0(shr_mem_16_cns_R1)
    );
  unreg_hier_69 unreg_34 (
      .in_0(shr_mem_17_cns_S0_iff),
      .out_0(shr_mem_17_cns_R0)
    );
  unreg_hier_69 unreg_35 (
      .in_0(shr_mem_17_cns_S1_iff),
      .out_0(shr_mem_17_cns_R1)
    );
  double_buffeaIgYu_0_cns_bctl double_buffeaIgYu_0_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(1'b0),
      .dout_0_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_0_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_0_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_0_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_0_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_0_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_0_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_0_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz),
      .din_0_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(1'b0),
      .din_0_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_0_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_0_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_0_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_0_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_0_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_0_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_0_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz),
      .din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .dout_0_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_0_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_0_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_0_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_1_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_1_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_2_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_2_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_3_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_3_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_4_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_4_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_5_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_5_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_6_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_6_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_7_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_7_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_8_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_8_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_9_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_9_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_10_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_10_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_11_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_11_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_12_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_12_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_13_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_13_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_14_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_14_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_15_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_15_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_16_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_16_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(1'b0),
      .dout_17_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(1'b0),
      .din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(1'b0),
      .din_17_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(1'b0),
      .dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_0_cns_S0(shr_mem_0_cns_S0_dmo),
      .shr_mem_0_cns_R0(shr_mem_0_cns_R0),
      .shr_mem_0_cns_S1(shr_mem_0_cns_S1_dmo),
      .shr_mem_0_cns_R1(shr_mem_0_cns_R1),
      .shr_mem_0_cns_addra_shi0(shr_mem_0_cns_addra_shi0),
      .shr_mem_0_cns_addra_shi1(shr_mem_0_cns_addra_shi1),
      .shr_mem_0_cns_addrb_shi0(shr_mem_0_cns_addrb_shi0),
      .shr_mem_0_cns_addrb_shi1(shr_mem_0_cns_addrb_shi1),
      .shr_mem_0_cns_csa_n_shi0(shr_mem_0_cns_csa_n_shi0),
      .shr_mem_0_cns_csa_n_shi1(shr_mem_0_cns_csa_n_shi1),
      .shr_mem_0_cns_csb_n_shi0(shr_mem_0_cns_csb_n_shi0),
      .shr_mem_0_cns_csb_n_shi1(shr_mem_0_cns_csb_n_shi1),
      .shr_mem_0_cns_dinb_shi0(shr_mem_0_cns_dinb_shi0),
      .shr_mem_0_cns_dinb_shi1(shr_mem_0_cns_dinb_shi1),
      .shr_mem_0_cns_douta_sho0(shr_mem_0_cns_douta_sho0),
      .shr_mem_0_cns_douta_sho1(shr_mem_0_cns_douta_sho1),
      .shr_mem_0_cns_S1_pff(shr_mem_0_cns_S1_iff),
      .shr_mem_0_cns_S0_pff(shr_mem_0_cns_S0_iff),
      .din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff)
    );
  double_buffeaIgYu_1_cns_bctl double_buffeaIgYu_1_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_1_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_1_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_1_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_1_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_1_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_1_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_1_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_1_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_1_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_1_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_1_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_1_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_1_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_1_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_1_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_1_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_1_cns_S0(shr_mem_1_cns_S0_dmo),
      .shr_mem_1_cns_R0(shr_mem_1_cns_R0),
      .shr_mem_1_cns_S1(shr_mem_1_cns_S1_dmo),
      .shr_mem_1_cns_R1(shr_mem_1_cns_R1),
      .shr_mem_1_cns_addra_shi0(shr_mem_1_cns_addra_shi0),
      .shr_mem_1_cns_addra_shi1(shr_mem_1_cns_addra_shi1),
      .shr_mem_1_cns_addrb_shi0(shr_mem_1_cns_addrb_shi0),
      .shr_mem_1_cns_addrb_shi1(shr_mem_1_cns_addrb_shi1),
      .shr_mem_1_cns_csa_n_shi0(shr_mem_1_cns_csa_n_shi0),
      .shr_mem_1_cns_csa_n_shi1(shr_mem_1_cns_csa_n_shi1),
      .shr_mem_1_cns_csb_n_shi0(shr_mem_1_cns_csb_n_shi0),
      .shr_mem_1_cns_csb_n_shi1(shr_mem_1_cns_csb_n_shi1),
      .shr_mem_1_cns_dinb_shi0(shr_mem_1_cns_dinb_shi0),
      .shr_mem_1_cns_dinb_shi1(shr_mem_1_cns_dinb_shi1),
      .shr_mem_1_cns_douta_sho0(shr_mem_1_cns_douta_sho0),
      .shr_mem_1_cns_douta_sho1(shr_mem_1_cns_douta_sho1),
      .shr_mem_1_cns_S1_pff(shr_mem_1_cns_S1_iff),
      .din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_1_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_1_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_1_cns_S0_pff(shr_mem_1_cns_S0_iff)
    );
  double_buffeaIgYu_2_cns_bctl double_buffeaIgYu_2_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_2_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_2_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_2_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_2_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_2_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_2_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_2_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_2_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_2_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_2_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_2_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_2_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_2_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_2_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_2_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_2_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_2_cns_S0(shr_mem_2_cns_S0_dmo),
      .shr_mem_2_cns_R0(shr_mem_2_cns_R0),
      .shr_mem_2_cns_S1(shr_mem_2_cns_S1_dmo),
      .shr_mem_2_cns_R1(shr_mem_2_cns_R1),
      .shr_mem_2_cns_addra_shi0(shr_mem_2_cns_addra_shi0),
      .shr_mem_2_cns_addra_shi1(shr_mem_2_cns_addra_shi1),
      .shr_mem_2_cns_addrb_shi0(shr_mem_2_cns_addrb_shi0),
      .shr_mem_2_cns_addrb_shi1(shr_mem_2_cns_addrb_shi1),
      .shr_mem_2_cns_csa_n_shi0(shr_mem_2_cns_csa_n_shi0),
      .shr_mem_2_cns_csa_n_shi1(shr_mem_2_cns_csa_n_shi1),
      .shr_mem_2_cns_csb_n_shi0(shr_mem_2_cns_csb_n_shi0),
      .shr_mem_2_cns_csb_n_shi1(shr_mem_2_cns_csb_n_shi1),
      .shr_mem_2_cns_dinb_shi0(shr_mem_2_cns_dinb_shi0),
      .shr_mem_2_cns_dinb_shi1(shr_mem_2_cns_dinb_shi1),
      .shr_mem_2_cns_douta_sho0(shr_mem_2_cns_douta_sho0),
      .shr_mem_2_cns_douta_sho1(shr_mem_2_cns_douta_sho1),
      .shr_mem_2_cns_S1_pff(shr_mem_2_cns_S1_iff),
      .din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_2_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_2_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_2_cns_S0_pff(shr_mem_2_cns_S0_iff)
    );
  double_buffeaIgYu_3_cns_bctl double_buffeaIgYu_3_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_3_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_3_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_3_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_3_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_3_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_3_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_3_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_3_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_3_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_3_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_3_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_3_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_3_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_3_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_3_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_3_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_3_cns_S0(shr_mem_3_cns_S0_dmo),
      .shr_mem_3_cns_R0(shr_mem_3_cns_R0),
      .shr_mem_3_cns_S1(shr_mem_3_cns_S1_dmo),
      .shr_mem_3_cns_R1(shr_mem_3_cns_R1),
      .shr_mem_3_cns_addra_shi0(shr_mem_3_cns_addra_shi0),
      .shr_mem_3_cns_addra_shi1(shr_mem_3_cns_addra_shi1),
      .shr_mem_3_cns_addrb_shi0(shr_mem_3_cns_addrb_shi0),
      .shr_mem_3_cns_addrb_shi1(shr_mem_3_cns_addrb_shi1),
      .shr_mem_3_cns_csa_n_shi0(shr_mem_3_cns_csa_n_shi0),
      .shr_mem_3_cns_csa_n_shi1(shr_mem_3_cns_csa_n_shi1),
      .shr_mem_3_cns_csb_n_shi0(shr_mem_3_cns_csb_n_shi0),
      .shr_mem_3_cns_csb_n_shi1(shr_mem_3_cns_csb_n_shi1),
      .shr_mem_3_cns_dinb_shi0(shr_mem_3_cns_dinb_shi0),
      .shr_mem_3_cns_dinb_shi1(shr_mem_3_cns_dinb_shi1),
      .shr_mem_3_cns_douta_sho0(shr_mem_3_cns_douta_sho0),
      .shr_mem_3_cns_douta_sho1(shr_mem_3_cns_douta_sho1),
      .shr_mem_3_cns_S1_pff(shr_mem_3_cns_S1_iff),
      .din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_3_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_3_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_3_cns_S0_pff(shr_mem_3_cns_S0_iff)
    );
  double_buffeaIgYu_4_cns_bctl double_buffeaIgYu_4_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_4_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_4_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_4_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_4_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_4_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_4_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_4_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_4_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_4_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_4_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_4_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_4_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_4_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_4_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_4_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_4_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_4_cns_S0(shr_mem_4_cns_S0_dmo),
      .shr_mem_4_cns_R0(shr_mem_4_cns_R0),
      .shr_mem_4_cns_S1(shr_mem_4_cns_S1_dmo),
      .shr_mem_4_cns_R1(shr_mem_4_cns_R1),
      .shr_mem_4_cns_addra_shi0(shr_mem_4_cns_addra_shi0),
      .shr_mem_4_cns_addra_shi1(shr_mem_4_cns_addra_shi1),
      .shr_mem_4_cns_addrb_shi0(shr_mem_4_cns_addrb_shi0),
      .shr_mem_4_cns_addrb_shi1(shr_mem_4_cns_addrb_shi1),
      .shr_mem_4_cns_csa_n_shi0(shr_mem_4_cns_csa_n_shi0),
      .shr_mem_4_cns_csa_n_shi1(shr_mem_4_cns_csa_n_shi1),
      .shr_mem_4_cns_csb_n_shi0(shr_mem_4_cns_csb_n_shi0),
      .shr_mem_4_cns_csb_n_shi1(shr_mem_4_cns_csb_n_shi1),
      .shr_mem_4_cns_dinb_shi0(shr_mem_4_cns_dinb_shi0),
      .shr_mem_4_cns_dinb_shi1(shr_mem_4_cns_dinb_shi1),
      .shr_mem_4_cns_douta_sho0(shr_mem_4_cns_douta_sho0),
      .shr_mem_4_cns_douta_sho1(shr_mem_4_cns_douta_sho1),
      .shr_mem_4_cns_S1_pff(shr_mem_4_cns_S1_iff),
      .din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_4_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_4_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_4_cns_S0_pff(shr_mem_4_cns_S0_iff)
    );
  double_buffeaIgYu_5_cns_bctl double_buffeaIgYu_5_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_5_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_5_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_5_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_5_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_5_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_5_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_5_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_5_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_5_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_5_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_5_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_5_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_5_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_5_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_5_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_5_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_5_cns_S0(shr_mem_5_cns_S0_dmo),
      .shr_mem_5_cns_R0(shr_mem_5_cns_R0),
      .shr_mem_5_cns_S1(shr_mem_5_cns_S1_dmo),
      .shr_mem_5_cns_R1(shr_mem_5_cns_R1),
      .shr_mem_5_cns_addra_shi0(shr_mem_5_cns_addra_shi0),
      .shr_mem_5_cns_addra_shi1(shr_mem_5_cns_addra_shi1),
      .shr_mem_5_cns_addrb_shi0(shr_mem_5_cns_addrb_shi0),
      .shr_mem_5_cns_addrb_shi1(shr_mem_5_cns_addrb_shi1),
      .shr_mem_5_cns_csa_n_shi0(shr_mem_5_cns_csa_n_shi0),
      .shr_mem_5_cns_csa_n_shi1(shr_mem_5_cns_csa_n_shi1),
      .shr_mem_5_cns_csb_n_shi0(shr_mem_5_cns_csb_n_shi0),
      .shr_mem_5_cns_csb_n_shi1(shr_mem_5_cns_csb_n_shi1),
      .shr_mem_5_cns_dinb_shi0(shr_mem_5_cns_dinb_shi0),
      .shr_mem_5_cns_dinb_shi1(shr_mem_5_cns_dinb_shi1),
      .shr_mem_5_cns_douta_sho0(shr_mem_5_cns_douta_sho0),
      .shr_mem_5_cns_douta_sho1(shr_mem_5_cns_douta_sho1),
      .shr_mem_5_cns_S1_pff(shr_mem_5_cns_S1_iff),
      .din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_5_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_5_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_5_cns_S0_pff(shr_mem_5_cns_S0_iff)
    );
  double_buffeaIgYu_6_cns_bctl double_buffeaIgYu_6_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_6_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_6_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_6_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_6_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_6_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_6_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_6_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_6_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_6_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_6_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_6_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_6_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_6_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_6_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_6_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_6_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_6_cns_S0(shr_mem_6_cns_S0_dmo),
      .shr_mem_6_cns_R0(shr_mem_6_cns_R0),
      .shr_mem_6_cns_S1(shr_mem_6_cns_S1_dmo),
      .shr_mem_6_cns_R1(shr_mem_6_cns_R1),
      .shr_mem_6_cns_addra_shi0(shr_mem_6_cns_addra_shi0),
      .shr_mem_6_cns_addra_shi1(shr_mem_6_cns_addra_shi1),
      .shr_mem_6_cns_addrb_shi0(shr_mem_6_cns_addrb_shi0),
      .shr_mem_6_cns_addrb_shi1(shr_mem_6_cns_addrb_shi1),
      .shr_mem_6_cns_csa_n_shi0(shr_mem_6_cns_csa_n_shi0),
      .shr_mem_6_cns_csa_n_shi1(shr_mem_6_cns_csa_n_shi1),
      .shr_mem_6_cns_csb_n_shi0(shr_mem_6_cns_csb_n_shi0),
      .shr_mem_6_cns_csb_n_shi1(shr_mem_6_cns_csb_n_shi1),
      .shr_mem_6_cns_dinb_shi0(shr_mem_6_cns_dinb_shi0),
      .shr_mem_6_cns_dinb_shi1(shr_mem_6_cns_dinb_shi1),
      .shr_mem_6_cns_douta_sho0(shr_mem_6_cns_douta_sho0),
      .shr_mem_6_cns_douta_sho1(shr_mem_6_cns_douta_sho1),
      .shr_mem_6_cns_S1_pff(shr_mem_6_cns_S1_iff),
      .din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_6_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_6_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_6_cns_S0_pff(shr_mem_6_cns_S0_iff)
    );
  double_buffeaIgYu_7_cns_bctl double_buffeaIgYu_7_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_7_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_7_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_7_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_7_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_7_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_7_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_7_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_7_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_7_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_7_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_7_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_7_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_7_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_7_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_7_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_7_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_7_cns_S0(shr_mem_7_cns_S0_dmo),
      .shr_mem_7_cns_R0(shr_mem_7_cns_R0),
      .shr_mem_7_cns_S1(shr_mem_7_cns_S1_dmo),
      .shr_mem_7_cns_R1(shr_mem_7_cns_R1),
      .shr_mem_7_cns_addra_shi0(shr_mem_7_cns_addra_shi0),
      .shr_mem_7_cns_addra_shi1(shr_mem_7_cns_addra_shi1),
      .shr_mem_7_cns_addrb_shi0(shr_mem_7_cns_addrb_shi0),
      .shr_mem_7_cns_addrb_shi1(shr_mem_7_cns_addrb_shi1),
      .shr_mem_7_cns_csa_n_shi0(shr_mem_7_cns_csa_n_shi0),
      .shr_mem_7_cns_csa_n_shi1(shr_mem_7_cns_csa_n_shi1),
      .shr_mem_7_cns_csb_n_shi0(shr_mem_7_cns_csb_n_shi0),
      .shr_mem_7_cns_csb_n_shi1(shr_mem_7_cns_csb_n_shi1),
      .shr_mem_7_cns_dinb_shi0(shr_mem_7_cns_dinb_shi0),
      .shr_mem_7_cns_dinb_shi1(shr_mem_7_cns_dinb_shi1),
      .shr_mem_7_cns_douta_sho0(shr_mem_7_cns_douta_sho0),
      .shr_mem_7_cns_douta_sho1(shr_mem_7_cns_douta_sho1),
      .shr_mem_7_cns_S1_pff(shr_mem_7_cns_S1_iff),
      .din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_7_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_7_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_7_cns_S0_pff(shr_mem_7_cns_S0_iff)
    );
  double_buffeaIgYu_8_cns_bctl double_buffeaIgYu_8_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_8_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_8_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_8_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_8_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_8_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_8_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_8_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_8_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_8_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_8_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_8_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_8_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_8_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_8_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_8_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_8_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_8_cns_S0(shr_mem_8_cns_S0_dmo),
      .shr_mem_8_cns_R0(shr_mem_8_cns_R0),
      .shr_mem_8_cns_S1(shr_mem_8_cns_S1_dmo),
      .shr_mem_8_cns_R1(shr_mem_8_cns_R1),
      .shr_mem_8_cns_addra_shi0(shr_mem_8_cns_addra_shi0),
      .shr_mem_8_cns_addra_shi1(shr_mem_8_cns_addra_shi1),
      .shr_mem_8_cns_addrb_shi0(shr_mem_8_cns_addrb_shi0),
      .shr_mem_8_cns_addrb_shi1(shr_mem_8_cns_addrb_shi1),
      .shr_mem_8_cns_csa_n_shi0(shr_mem_8_cns_csa_n_shi0),
      .shr_mem_8_cns_csa_n_shi1(shr_mem_8_cns_csa_n_shi1),
      .shr_mem_8_cns_csb_n_shi0(shr_mem_8_cns_csb_n_shi0),
      .shr_mem_8_cns_csb_n_shi1(shr_mem_8_cns_csb_n_shi1),
      .shr_mem_8_cns_dinb_shi0(shr_mem_8_cns_dinb_shi0),
      .shr_mem_8_cns_dinb_shi1(shr_mem_8_cns_dinb_shi1),
      .shr_mem_8_cns_douta_sho0(shr_mem_8_cns_douta_sho0),
      .shr_mem_8_cns_douta_sho1(shr_mem_8_cns_douta_sho1),
      .shr_mem_8_cns_S1_pff(shr_mem_8_cns_S1_iff),
      .din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_8_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_8_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_8_cns_S0_pff(shr_mem_8_cns_S0_iff)
    );
  double_buffeaIgYu_9_cns_bctl double_buffeaIgYu_9_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_9_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_9_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_9_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_9_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_9_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_9_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_9_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_9_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_9_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_9_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_9_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_9_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_9_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_9_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_9_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_9_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_9_cns_S0(shr_mem_9_cns_S0_dmo),
      .shr_mem_9_cns_R0(shr_mem_9_cns_R0),
      .shr_mem_9_cns_S1(shr_mem_9_cns_S1_dmo),
      .shr_mem_9_cns_R1(shr_mem_9_cns_R1),
      .shr_mem_9_cns_addra_shi0(shr_mem_9_cns_addra_shi0),
      .shr_mem_9_cns_addra_shi1(shr_mem_9_cns_addra_shi1),
      .shr_mem_9_cns_addrb_shi0(shr_mem_9_cns_addrb_shi0),
      .shr_mem_9_cns_addrb_shi1(shr_mem_9_cns_addrb_shi1),
      .shr_mem_9_cns_csa_n_shi0(shr_mem_9_cns_csa_n_shi0),
      .shr_mem_9_cns_csa_n_shi1(shr_mem_9_cns_csa_n_shi1),
      .shr_mem_9_cns_csb_n_shi0(shr_mem_9_cns_csb_n_shi0),
      .shr_mem_9_cns_csb_n_shi1(shr_mem_9_cns_csb_n_shi1),
      .shr_mem_9_cns_dinb_shi0(shr_mem_9_cns_dinb_shi0),
      .shr_mem_9_cns_dinb_shi1(shr_mem_9_cns_dinb_shi1),
      .shr_mem_9_cns_douta_sho0(shr_mem_9_cns_douta_sho0),
      .shr_mem_9_cns_douta_sho1(shr_mem_9_cns_douta_sho1),
      .shr_mem_9_cns_S1_pff(shr_mem_9_cns_S1_iff),
      .din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_9_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_9_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_9_cns_S0_pff(shr_mem_9_cns_S0_iff)
    );
  double_buffeoFsRV10_cns_bctl double_buffeoFsRV10_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_10_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_10_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_10_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_10_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_10_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_10_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_10_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_10_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_10_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_10_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_10_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_10_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_10_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_10_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_10_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_10_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_10_cns_S0(shr_mem_10_cns_S0_dmo),
      .shr_mem_10_cns_R0(shr_mem_10_cns_R0),
      .shr_mem_10_cns_S1(shr_mem_10_cns_S1_dmo),
      .shr_mem_10_cns_R1(shr_mem_10_cns_R1),
      .shr_mem_10_cns_addra_shi0(shr_mem_10_cns_addra_shi0),
      .shr_mem_10_cns_addra_shi1(shr_mem_10_cns_addra_shi1),
      .shr_mem_10_cns_addrb_shi0(shr_mem_10_cns_addrb_shi0),
      .shr_mem_10_cns_addrb_shi1(shr_mem_10_cns_addrb_shi1),
      .shr_mem_10_cns_csa_n_shi0(shr_mem_10_cns_csa_n_shi0),
      .shr_mem_10_cns_csa_n_shi1(shr_mem_10_cns_csa_n_shi1),
      .shr_mem_10_cns_csb_n_shi0(shr_mem_10_cns_csb_n_shi0),
      .shr_mem_10_cns_csb_n_shi1(shr_mem_10_cns_csb_n_shi1),
      .shr_mem_10_cns_dinb_shi0(shr_mem_10_cns_dinb_shi0),
      .shr_mem_10_cns_dinb_shi1(shr_mem_10_cns_dinb_shi1),
      .shr_mem_10_cns_douta_sho0(shr_mem_10_cns_douta_sho0),
      .shr_mem_10_cns_douta_sho1(shr_mem_10_cns_douta_sho1),
      .shr_mem_10_cns_S1_pff(shr_mem_10_cns_S1_iff),
      .din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_10_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_10_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_10_cns_S0_pff(shr_mem_10_cns_S0_iff)
    );
  double_buffeoFsRV11_cns_bctl double_buffeoFsRV11_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_11_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_11_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_11_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_11_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_11_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_11_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_11_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_11_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_11_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_11_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_11_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_11_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_11_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_11_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_11_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_11_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_11_cns_S0(shr_mem_11_cns_S0_dmo),
      .shr_mem_11_cns_R0(shr_mem_11_cns_R0),
      .shr_mem_11_cns_S1(shr_mem_11_cns_S1_dmo),
      .shr_mem_11_cns_R1(shr_mem_11_cns_R1),
      .shr_mem_11_cns_addra_shi0(shr_mem_11_cns_addra_shi0),
      .shr_mem_11_cns_addra_shi1(shr_mem_11_cns_addra_shi1),
      .shr_mem_11_cns_addrb_shi0(shr_mem_11_cns_addrb_shi0),
      .shr_mem_11_cns_addrb_shi1(shr_mem_11_cns_addrb_shi1),
      .shr_mem_11_cns_csa_n_shi0(shr_mem_11_cns_csa_n_shi0),
      .shr_mem_11_cns_csa_n_shi1(shr_mem_11_cns_csa_n_shi1),
      .shr_mem_11_cns_csb_n_shi0(shr_mem_11_cns_csb_n_shi0),
      .shr_mem_11_cns_csb_n_shi1(shr_mem_11_cns_csb_n_shi1),
      .shr_mem_11_cns_dinb_shi0(shr_mem_11_cns_dinb_shi0),
      .shr_mem_11_cns_dinb_shi1(shr_mem_11_cns_dinb_shi1),
      .shr_mem_11_cns_douta_sho0(shr_mem_11_cns_douta_sho0),
      .shr_mem_11_cns_douta_sho1(shr_mem_11_cns_douta_sho1),
      .shr_mem_11_cns_S1_pff(shr_mem_11_cns_S1_iff),
      .din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_11_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_11_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_11_cns_S0_pff(shr_mem_11_cns_S0_iff)
    );
  double_buffeoFsRV12_cns_bctl double_buffeoFsRV12_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_12_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_12_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_12_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_12_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_12_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_12_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_12_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_12_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_12_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_12_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_12_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_12_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_12_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_12_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_12_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_12_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_12_cns_S0(shr_mem_12_cns_S0_dmo),
      .shr_mem_12_cns_R0(shr_mem_12_cns_R0),
      .shr_mem_12_cns_S1(shr_mem_12_cns_S1_dmo),
      .shr_mem_12_cns_R1(shr_mem_12_cns_R1),
      .shr_mem_12_cns_addra_shi0(shr_mem_12_cns_addra_shi0),
      .shr_mem_12_cns_addra_shi1(shr_mem_12_cns_addra_shi1),
      .shr_mem_12_cns_addrb_shi0(shr_mem_12_cns_addrb_shi0),
      .shr_mem_12_cns_addrb_shi1(shr_mem_12_cns_addrb_shi1),
      .shr_mem_12_cns_csa_n_shi0(shr_mem_12_cns_csa_n_shi0),
      .shr_mem_12_cns_csa_n_shi1(shr_mem_12_cns_csa_n_shi1),
      .shr_mem_12_cns_csb_n_shi0(shr_mem_12_cns_csb_n_shi0),
      .shr_mem_12_cns_csb_n_shi1(shr_mem_12_cns_csb_n_shi1),
      .shr_mem_12_cns_dinb_shi0(shr_mem_12_cns_dinb_shi0),
      .shr_mem_12_cns_dinb_shi1(shr_mem_12_cns_dinb_shi1),
      .shr_mem_12_cns_douta_sho0(shr_mem_12_cns_douta_sho0),
      .shr_mem_12_cns_douta_sho1(shr_mem_12_cns_douta_sho1),
      .shr_mem_12_cns_S1_pff(shr_mem_12_cns_S1_iff),
      .din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_12_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_12_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_12_cns_S0_pff(shr_mem_12_cns_S0_iff)
    );
  double_buffeoFsRV13_cns_bctl double_buffeoFsRV13_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_13_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_13_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_13_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_13_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_13_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_13_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_13_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_13_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_13_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_13_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_13_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_13_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_13_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_13_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_13_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_13_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_13_cns_S0(shr_mem_13_cns_S0_dmo),
      .shr_mem_13_cns_R0(shr_mem_13_cns_R0),
      .shr_mem_13_cns_S1(shr_mem_13_cns_S1_dmo),
      .shr_mem_13_cns_R1(shr_mem_13_cns_R1),
      .shr_mem_13_cns_addra_shi0(shr_mem_13_cns_addra_shi0),
      .shr_mem_13_cns_addra_shi1(shr_mem_13_cns_addra_shi1),
      .shr_mem_13_cns_addrb_shi0(shr_mem_13_cns_addrb_shi0),
      .shr_mem_13_cns_addrb_shi1(shr_mem_13_cns_addrb_shi1),
      .shr_mem_13_cns_csa_n_shi0(shr_mem_13_cns_csa_n_shi0),
      .shr_mem_13_cns_csa_n_shi1(shr_mem_13_cns_csa_n_shi1),
      .shr_mem_13_cns_csb_n_shi0(shr_mem_13_cns_csb_n_shi0),
      .shr_mem_13_cns_csb_n_shi1(shr_mem_13_cns_csb_n_shi1),
      .shr_mem_13_cns_dinb_shi0(shr_mem_13_cns_dinb_shi0),
      .shr_mem_13_cns_dinb_shi1(shr_mem_13_cns_dinb_shi1),
      .shr_mem_13_cns_douta_sho0(shr_mem_13_cns_douta_sho0),
      .shr_mem_13_cns_douta_sho1(shr_mem_13_cns_douta_sho1),
      .shr_mem_13_cns_S1_pff(shr_mem_13_cns_S1_iff),
      .din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_13_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_13_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_13_cns_S0_pff(shr_mem_13_cns_S0_iff)
    );
  double_buffeoFsRV14_cns_bctl double_buffeoFsRV14_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_14_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_14_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_14_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_14_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_14_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_14_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_14_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_14_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_14_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_14_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_14_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_14_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_14_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_14_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_14_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_14_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_14_cns_S0(shr_mem_14_cns_S0_dmo),
      .shr_mem_14_cns_R0(shr_mem_14_cns_R0),
      .shr_mem_14_cns_S1(shr_mem_14_cns_S1_dmo),
      .shr_mem_14_cns_R1(shr_mem_14_cns_R1),
      .shr_mem_14_cns_addra_shi0(shr_mem_14_cns_addra_shi0),
      .shr_mem_14_cns_addra_shi1(shr_mem_14_cns_addra_shi1),
      .shr_mem_14_cns_addrb_shi0(shr_mem_14_cns_addrb_shi0),
      .shr_mem_14_cns_addrb_shi1(shr_mem_14_cns_addrb_shi1),
      .shr_mem_14_cns_csa_n_shi0(shr_mem_14_cns_csa_n_shi0),
      .shr_mem_14_cns_csa_n_shi1(shr_mem_14_cns_csa_n_shi1),
      .shr_mem_14_cns_csb_n_shi0(shr_mem_14_cns_csb_n_shi0),
      .shr_mem_14_cns_csb_n_shi1(shr_mem_14_cns_csb_n_shi1),
      .shr_mem_14_cns_dinb_shi0(shr_mem_14_cns_dinb_shi0),
      .shr_mem_14_cns_dinb_shi1(shr_mem_14_cns_dinb_shi1),
      .shr_mem_14_cns_douta_sho0(shr_mem_14_cns_douta_sho0),
      .shr_mem_14_cns_douta_sho1(shr_mem_14_cns_douta_sho1),
      .shr_mem_14_cns_S1_pff(shr_mem_14_cns_S1_iff),
      .din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_14_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_14_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_14_cns_S0_pff(shr_mem_14_cns_S0_iff)
    );
  double_buffeoFsRV15_cns_bctl double_buffeoFsRV15_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_15_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_15_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_15_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_15_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_15_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_15_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_15_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_15_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_15_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_15_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_15_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_15_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_15_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_15_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_15_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_15_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_15_cns_S0(shr_mem_15_cns_S0_dmo),
      .shr_mem_15_cns_R0(shr_mem_15_cns_R0),
      .shr_mem_15_cns_S1(shr_mem_15_cns_S1_dmo),
      .shr_mem_15_cns_R1(shr_mem_15_cns_R1),
      .shr_mem_15_cns_addra_shi0(shr_mem_15_cns_addra_shi0),
      .shr_mem_15_cns_addra_shi1(shr_mem_15_cns_addra_shi1),
      .shr_mem_15_cns_addrb_shi0(shr_mem_15_cns_addrb_shi0),
      .shr_mem_15_cns_addrb_shi1(shr_mem_15_cns_addrb_shi1),
      .shr_mem_15_cns_csa_n_shi0(shr_mem_15_cns_csa_n_shi0),
      .shr_mem_15_cns_csa_n_shi1(shr_mem_15_cns_csa_n_shi1),
      .shr_mem_15_cns_csb_n_shi0(shr_mem_15_cns_csb_n_shi0),
      .shr_mem_15_cns_csb_n_shi1(shr_mem_15_cns_csb_n_shi1),
      .shr_mem_15_cns_dinb_shi0(shr_mem_15_cns_dinb_shi0),
      .shr_mem_15_cns_dinb_shi1(shr_mem_15_cns_dinb_shi1),
      .shr_mem_15_cns_douta_sho0(shr_mem_15_cns_douta_sho0),
      .shr_mem_15_cns_douta_sho1(shr_mem_15_cns_douta_sho1),
      .shr_mem_15_cns_S1_pff(shr_mem_15_cns_S1_iff),
      .din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_15_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_15_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_15_cns_S0_pff(shr_mem_15_cns_S0_iff)
    );
  double_buffeoFsRV16_cns_bctl double_buffeoFsRV16_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_16_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_16_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_16_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_16_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_16_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_16_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_16_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_16_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_16_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_16_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_16_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_16_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_16_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_16_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_16_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_16_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_16_cns_S0(shr_mem_16_cns_S0_dmo),
      .shr_mem_16_cns_R0(shr_mem_16_cns_R0),
      .shr_mem_16_cns_S1(shr_mem_16_cns_S1_dmo),
      .shr_mem_16_cns_R1(shr_mem_16_cns_R1),
      .shr_mem_16_cns_addra_shi0(shr_mem_16_cns_addra_shi0),
      .shr_mem_16_cns_addra_shi1(shr_mem_16_cns_addra_shi1),
      .shr_mem_16_cns_addrb_shi0(shr_mem_16_cns_addrb_shi0),
      .shr_mem_16_cns_addrb_shi1(shr_mem_16_cns_addrb_shi1),
      .shr_mem_16_cns_csa_n_shi0(shr_mem_16_cns_csa_n_shi0),
      .shr_mem_16_cns_csa_n_shi1(shr_mem_16_cns_csa_n_shi1),
      .shr_mem_16_cns_csb_n_shi0(shr_mem_16_cns_csb_n_shi0),
      .shr_mem_16_cns_csb_n_shi1(shr_mem_16_cns_csb_n_shi1),
      .shr_mem_16_cns_dinb_shi0(shr_mem_16_cns_dinb_shi0),
      .shr_mem_16_cns_dinb_shi1(shr_mem_16_cns_dinb_shi1),
      .shr_mem_16_cns_douta_sho0(shr_mem_16_cns_douta_sho0),
      .shr_mem_16_cns_douta_sho1(shr_mem_16_cns_douta_sho1),
      .shr_mem_16_cns_S1_pff(shr_mem_16_cns_S1_iff),
      .din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_16_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_16_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_16_cns_S0_pff(shr_mem_16_cns_S0_iff)
    );
  double_buffeoFsRV17_cns_bctl double_buffeoFsRV17_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_addra_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(7'b0),
      .dout_17_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_17_rsc_addrb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_17_rsc_dinb_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_17_rsc_douta_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst(dout_17_rsc_req_vz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst),
      .dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz(1'b0),
      .din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_addra_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(7'b0),
      .din_17_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_17_rsc_addrb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_17_rsc_dinb_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_17_rsc_douta_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst(din_17_rsc_req_vz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst),
      .din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz(1'b0),
      .dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud(dout_17_rsc_csa_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud),
      .dout_17_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud(dout_17_rsc_rls_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_bud),
      .din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud(din_17_rsc_csa_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud),
      .din_17_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud(din_17_rsc_rls_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_bud),
      .shr_mem_17_cns_S0(shr_mem_17_cns_S0_dmo),
      .shr_mem_17_cns_R0(shr_mem_17_cns_R0),
      .shr_mem_17_cns_S1(shr_mem_17_cns_S1_dmo),
      .shr_mem_17_cns_R1(shr_mem_17_cns_R1),
      .shr_mem_17_cns_addra_shi0(shr_mem_17_cns_addra_shi0),
      .shr_mem_17_cns_addra_shi1(shr_mem_17_cns_addra_shi1),
      .shr_mem_17_cns_addrb_shi0(shr_mem_17_cns_addrb_shi0),
      .shr_mem_17_cns_addrb_shi1(shr_mem_17_cns_addrb_shi1),
      .shr_mem_17_cns_csa_n_shi0(shr_mem_17_cns_csa_n_shi0),
      .shr_mem_17_cns_csa_n_shi1(shr_mem_17_cns_csa_n_shi1),
      .shr_mem_17_cns_csb_n_shi0(shr_mem_17_cns_csb_n_shi0),
      .shr_mem_17_cns_csb_n_shi1(shr_mem_17_cns_csb_n_shi1),
      .shr_mem_17_cns_dinb_shi0(shr_mem_17_cns_dinb_shi0),
      .shr_mem_17_cns_dinb_shi1(shr_mem_17_cns_dinb_shi1),
      .shr_mem_17_cns_douta_sho0(shr_mem_17_cns_douta_sho0),
      .shr_mem_17_cns_douta_sho1(shr_mem_17_cns_douta_sho1),
      .shr_mem_17_cns_S1_pff(shr_mem_17_cns_S1_iff),
      .din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_pff(din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_iff),
      .din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_pff(din_17_rsc_csb_n_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst_buz_bud_iff),
      .dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_pff(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_iff),
      .dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_pff(dout_17_rsc_csb_n_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst_buz_bud_iff),
      .shr_mem_17_cns_S0_pff(shr_mem_17_cns_S0_iff)
    );
  assign din_rsc_lz = din_rsc_lz_nWRITE_BLOCK_INPUT_DTYPE_64_16_1_3_inst;
  assign dout_rsc_lz = dout_rsc_lz_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
  assign dout_rsc_z = dout_rsc_z_nREAD_BLOCK_INPUT_DTYPE_64_16_4_1_3_inst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffer_weights_DTYPE_2_16_4_1_3
// ------------------------------------------------------------------


module double_buffer_weights_DTYPE_2_16_4_1_3 (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, dout_rsc_z, dout_rsc_vz, dout_rsc_lz,
      clamp_mem, scan_n, shift_n, slp_nret_n, slp_ret_n
);
  input clk;
  input rst;
  input [63:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  output [63:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;
  input clamp_mem;
  input scan_n;
  input shift_n;
  input slp_nret_n;
  input slp_ret_n;


  // Interconnect Declarations
  wire din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  wire dout_rsc_csa_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  wire dout_rsc_csb_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  wire [6:0] dout_rsc_addra_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  wire [6:0] dout_rsc_addrb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  wire [63:0] dout_rsc_dinb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  wire [63:0] dout_rsc_douta_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  wire dout_rsc_req_vz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  wire din_rsc_csa_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  wire din_rsc_csb_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  wire [6:0] din_rsc_addra_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  wire [6:0] din_rsc_addrb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  wire [63:0] din_rsc_dinb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  wire [63:0] din_rsc_douta_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  wire din_rsc_req_vz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  wire [63:0] dout_rsc_z_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  wire dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  wire din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud;
  wire dout_rsc_rls_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud;
  wire din_rsc_rls_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud;
  wire dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud;
  wire shr_mem_cns_R0;
  wire shr_mem_cns_R1;
  wire [6:0] shr_mem_cns_addra_shi0;
  wire [6:0] shr_mem_cns_addra_shi1;
  wire [6:0] shr_mem_cns_addrb_shi0;
  wire [6:0] shr_mem_cns_addrb_shi1;
  wire shr_mem_cns_csa_n_shi0;
  wire shr_mem_cns_csa_n_shi1;
  wire shr_mem_cns_csb_n_shi0;
  wire shr_mem_cns_csb_n_shi1;
  wire [63:0] shr_mem_cns_dinb_shi0;
  wire [63:0] shr_mem_cns_dinb_shi1;
  wire [63:0] shr_mem_cns_douta_sho0;
  wire [63:0] shr_mem_cns_douta_sho1;
  wire shr_mem_cns_unc_1;
  wire shr_mem_cns_S1_iff;
  wire shr_mem_cns_S0_iff;
  wire shr_mem_cns_S0_dmo;
  wire shr_mem_cns_S1_dmo;


  // Interconnect Declarations for Component Instantiations 
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_cns_comp (
      .addra(shr_mem_cns_addra_shi0),
      .addrb(shr_mem_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_cns_csa_n_shi0),
      .csb_n(shr_mem_cns_csb_n_shi0),
      .dinb(shr_mem_cns_dinb_shi0),
      .douta(shr_mem_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_cns_unc_1)
    );
  cat_ram2p_half_128x64 #(.filename(-1073740000),
  .filename_size(32'sd0),
  .VLOG_DELAY(32'sd0),
  .MEMORY_ACC_WIDTH(32'sd0)) shr_mem_cns_comp_1 (
      .addra(shr_mem_cns_addra_shi1),
      .addrb(shr_mem_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_cns_csa_n_shi1),
      .csb_n(shr_mem_cns_csb_n_shi1),
      .dinb(shr_mem_cns_dinb_shi1),
      .douta(shr_mem_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_cns_unc_1)
    );
  WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_1 WRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(din_rsc_z),
      .din_rsc_vz(din_rsc_vz),
      .din_rsc_lz(din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud),
      .dout_rsc_csa_n(dout_rsc_csa_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_csb_n(dout_rsc_csb_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_addra(dout_rsc_addra_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_addrb(dout_rsc_addrb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_dinb(dout_rsc_dinb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_douta(dout_rsc_douta_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_req_vz(dout_rsc_req_vz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_rls_lz(dout_rsc_rls_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud)
    );
  READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_1 READ_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_csa_n(din_rsc_csa_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_csb_n(din_rsc_csb_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_addra(din_rsc_addra_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_addrb(din_rsc_addrb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_dinb(din_rsc_dinb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_douta(din_rsc_douta_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_req_vz(din_rsc_req_vz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_rls_lz(din_rsc_rls_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud),
      .dout_rsc_z(dout_rsc_z_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .dout_rsc_vz(dout_rsc_vz),
      .dout_rsc_lz(dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud)
    );
  unreg_hier_33 unreg (
      .in_0(shr_mem_cns_S0_iff),
      .out_0(shr_mem_cns_R0)
    );
  unreg_hier_33 unreg_1 (
      .in_0(shr_mem_cns_S1_iff),
      .out_0(shr_mem_cns_R1)
    );
  double_buffepBGdfem_cns_bctl double_buffepBGdfem_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst(din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_csa_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst(1'b0),
      .dout_rsc_csb_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst(dout_rsc_csb_n_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_addra_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst(7'b0),
      .dout_rsc_addrb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst(dout_rsc_addrb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_dinb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst(dout_rsc_dinb_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_douta_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst(dout_rsc_douta_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .dout_rsc_req_vz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst(dout_rsc_req_vz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst),
      .din_rsc_csa_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst(1'b0),
      .din_rsc_csb_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst(din_rsc_csb_n_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_addra_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst(7'b0),
      .din_rsc_addrb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst(din_rsc_addrb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_dinb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst(din_rsc_dinb_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_douta_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst(din_rsc_douta_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_req_vz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst(din_rsc_req_vz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst(dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst),
      .din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud(din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud),
      .dout_rsc_rls_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud(dout_rsc_rls_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst_bud),
      .din_rsc_rls_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud(din_rsc_rls_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud),
      .dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud(dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst_bud),
      .shr_mem_cns_S0(shr_mem_cns_S0_dmo),
      .shr_mem_cns_R0(shr_mem_cns_R0),
      .shr_mem_cns_S1(shr_mem_cns_S1_dmo),
      .shr_mem_cns_R1(shr_mem_cns_R1),
      .shr_mem_cns_addra_shi0(shr_mem_cns_addra_shi0),
      .shr_mem_cns_addra_shi1(shr_mem_cns_addra_shi1),
      .shr_mem_cns_addrb_shi0(shr_mem_cns_addrb_shi0),
      .shr_mem_cns_addrb_shi1(shr_mem_cns_addrb_shi1),
      .shr_mem_cns_csa_n_shi0(shr_mem_cns_csa_n_shi0),
      .shr_mem_cns_csa_n_shi1(shr_mem_cns_csa_n_shi1),
      .shr_mem_cns_csb_n_shi0(shr_mem_cns_csb_n_shi0),
      .shr_mem_cns_csb_n_shi1(shr_mem_cns_csb_n_shi1),
      .shr_mem_cns_dinb_shi0(shr_mem_cns_dinb_shi0),
      .shr_mem_cns_dinb_shi1(shr_mem_cns_dinb_shi1),
      .shr_mem_cns_douta_sho0(shr_mem_cns_douta_sho0),
      .shr_mem_cns_douta_sho1(shr_mem_cns_douta_sho1),
      .shr_mem_cns_S1_pff(shr_mem_cns_S1_iff),
      .shr_mem_cns_S0_pff(shr_mem_cns_S0_iff)
    );
  assign din_rsc_lz = din_rsc_lz_nWRITE_BLOCK_WEIGHTS_DTYPE_4_1_3_2_inst;
  assign dout_rsc_lz = dout_rsc_lz_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
  assign dout_rsc_z = dout_rsc_z_nREAD_BLOCK_WEIGHTS_DTYPE_16_4_1_3_2_inst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    double_buffer_output_DTYPE_2_16_64_4
// ------------------------------------------------------------------


module double_buffer_output_DTYPE_2_16_64_4 (
  clk, rst, din_rsc_z, din_rsc_vz, din_rsc_lz, dout_rsc_z, dout_rsc_vz, dout_rsc_lz,
      clamp_mem, scan_n, shift_n, slp_nret_n, slp_ret_n
);
  input clk;
  input rst;
  input [1023:0] din_rsc_z;
  input din_rsc_vz;
  output din_rsc_lz;
  output [1023:0] dout_rsc_z;
  input dout_rsc_vz;
  output dout_rsc_lz;
  input clamp_mem;
  input scan_n;
  input shift_n;
  input slp_nret_n;
  input slp_ret_n;


  // Interconnect Declarations
  wire din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_0_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_0_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_0_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_0_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_0_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_0_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_0_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_1_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_1_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_1_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_1_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_1_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_2_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_2_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_2_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_2_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_2_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_3_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_3_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_3_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_3_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_3_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_4_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_4_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_4_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_4_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_4_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_5_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_5_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_5_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_5_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_5_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_6_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_6_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_6_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_6_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_6_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_7_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_7_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_7_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_7_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_7_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_8_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_8_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_8_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_8_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_8_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_9_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_9_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_9_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_9_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_9_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_10_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_10_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_10_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_10_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_10_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_11_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_11_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_11_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_11_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_11_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_12_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_12_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_12_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_12_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_12_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_13_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_13_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_13_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_13_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_13_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_14_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_14_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_14_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_14_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_14_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_15_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] dout_15_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_15_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] dout_15_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_15_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_0_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_0_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_0_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_0_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_0_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_0_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_0_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_1_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_1_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_1_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_1_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_1_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_2_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_2_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_2_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_2_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_2_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_3_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_3_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_3_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_3_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_3_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_4_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_4_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_4_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_4_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_4_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_5_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_5_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_5_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_5_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_5_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_6_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_6_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_6_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_6_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_6_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_7_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_7_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_7_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_7_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_7_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_8_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_8_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_8_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_8_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_8_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_9_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_9_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_9_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_9_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_9_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_10_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_10_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_10_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_10_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_10_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_11_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_11_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_11_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_11_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_11_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_12_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_12_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_12_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_12_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_12_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_13_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_13_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_13_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_13_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_13_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_14_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_14_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_14_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_14_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_14_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_15_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [7:0] din_15_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_15_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [63:0] din_15_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_15_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire [1023:0] dout_rsc_z_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  wire din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz;
  wire din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_0_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_0_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_1_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_1_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_2_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_2_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_3_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_3_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_4_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_4_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_5_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_5_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_6_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_6_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_7_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_7_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_8_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_8_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_9_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_9_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_10_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_10_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_11_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_11_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_12_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_12_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_13_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_13_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_14_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_14_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire dout_15_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud;
  wire din_15_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud;
  wire shr_mem_0_cns_R0;
  wire shr_mem_0_cns_R1;
  wire [7:0] shr_mem_0_cns_addra_shi0;
  wire [7:0] shr_mem_0_cns_addra_shi1;
  wire [7:0] shr_mem_0_cns_addrb_shi0;
  wire [7:0] shr_mem_0_cns_addrb_shi1;
  wire shr_mem_0_cns_csa_n_shi0;
  wire shr_mem_0_cns_csa_n_shi1;
  wire shr_mem_0_cns_csb_n_shi0;
  wire shr_mem_0_cns_csb_n_shi1;
  wire [63:0] shr_mem_0_cns_dinb_shi0;
  wire [63:0] shr_mem_0_cns_dinb_shi1;
  wire [63:0] shr_mem_0_cns_douta_sho0;
  wire [63:0] shr_mem_0_cns_douta_sho1;
  wire shr_mem_0_cns_unc_1;
  wire shr_mem_1_cns_R0;
  wire shr_mem_1_cns_R1;
  wire [7:0] shr_mem_1_cns_addra_shi0;
  wire [7:0] shr_mem_1_cns_addra_shi1;
  wire [7:0] shr_mem_1_cns_addrb_shi0;
  wire [7:0] shr_mem_1_cns_addrb_shi1;
  wire shr_mem_1_cns_csa_n_shi0;
  wire shr_mem_1_cns_csa_n_shi1;
  wire shr_mem_1_cns_csb_n_shi0;
  wire shr_mem_1_cns_csb_n_shi1;
  wire [63:0] shr_mem_1_cns_dinb_shi0;
  wire [63:0] shr_mem_1_cns_dinb_shi1;
  wire [63:0] shr_mem_1_cns_douta_sho0;
  wire [63:0] shr_mem_1_cns_douta_sho1;
  wire shr_mem_1_cns_unc_1;
  wire shr_mem_2_cns_R0;
  wire shr_mem_2_cns_R1;
  wire [7:0] shr_mem_2_cns_addra_shi0;
  wire [7:0] shr_mem_2_cns_addra_shi1;
  wire [7:0] shr_mem_2_cns_addrb_shi0;
  wire [7:0] shr_mem_2_cns_addrb_shi1;
  wire shr_mem_2_cns_csa_n_shi0;
  wire shr_mem_2_cns_csa_n_shi1;
  wire shr_mem_2_cns_csb_n_shi0;
  wire shr_mem_2_cns_csb_n_shi1;
  wire [63:0] shr_mem_2_cns_dinb_shi0;
  wire [63:0] shr_mem_2_cns_dinb_shi1;
  wire [63:0] shr_mem_2_cns_douta_sho0;
  wire [63:0] shr_mem_2_cns_douta_sho1;
  wire shr_mem_2_cns_unc_1;
  wire shr_mem_3_cns_R0;
  wire shr_mem_3_cns_R1;
  wire [7:0] shr_mem_3_cns_addra_shi0;
  wire [7:0] shr_mem_3_cns_addra_shi1;
  wire [7:0] shr_mem_3_cns_addrb_shi0;
  wire [7:0] shr_mem_3_cns_addrb_shi1;
  wire shr_mem_3_cns_csa_n_shi0;
  wire shr_mem_3_cns_csa_n_shi1;
  wire shr_mem_3_cns_csb_n_shi0;
  wire shr_mem_3_cns_csb_n_shi1;
  wire [63:0] shr_mem_3_cns_dinb_shi0;
  wire [63:0] shr_mem_3_cns_dinb_shi1;
  wire [63:0] shr_mem_3_cns_douta_sho0;
  wire [63:0] shr_mem_3_cns_douta_sho1;
  wire shr_mem_3_cns_unc_1;
  wire shr_mem_4_cns_R0;
  wire shr_mem_4_cns_R1;
  wire [7:0] shr_mem_4_cns_addra_shi0;
  wire [7:0] shr_mem_4_cns_addra_shi1;
  wire [7:0] shr_mem_4_cns_addrb_shi0;
  wire [7:0] shr_mem_4_cns_addrb_shi1;
  wire shr_mem_4_cns_csa_n_shi0;
  wire shr_mem_4_cns_csa_n_shi1;
  wire shr_mem_4_cns_csb_n_shi0;
  wire shr_mem_4_cns_csb_n_shi1;
  wire [63:0] shr_mem_4_cns_dinb_shi0;
  wire [63:0] shr_mem_4_cns_dinb_shi1;
  wire [63:0] shr_mem_4_cns_douta_sho0;
  wire [63:0] shr_mem_4_cns_douta_sho1;
  wire shr_mem_4_cns_unc_1;
  wire shr_mem_5_cns_R0;
  wire shr_mem_5_cns_R1;
  wire [7:0] shr_mem_5_cns_addra_shi0;
  wire [7:0] shr_mem_5_cns_addra_shi1;
  wire [7:0] shr_mem_5_cns_addrb_shi0;
  wire [7:0] shr_mem_5_cns_addrb_shi1;
  wire shr_mem_5_cns_csa_n_shi0;
  wire shr_mem_5_cns_csa_n_shi1;
  wire shr_mem_5_cns_csb_n_shi0;
  wire shr_mem_5_cns_csb_n_shi1;
  wire [63:0] shr_mem_5_cns_dinb_shi0;
  wire [63:0] shr_mem_5_cns_dinb_shi1;
  wire [63:0] shr_mem_5_cns_douta_sho0;
  wire [63:0] shr_mem_5_cns_douta_sho1;
  wire shr_mem_5_cns_unc_1;
  wire shr_mem_6_cns_R0;
  wire shr_mem_6_cns_R1;
  wire [7:0] shr_mem_6_cns_addra_shi0;
  wire [7:0] shr_mem_6_cns_addra_shi1;
  wire [7:0] shr_mem_6_cns_addrb_shi0;
  wire [7:0] shr_mem_6_cns_addrb_shi1;
  wire shr_mem_6_cns_csa_n_shi0;
  wire shr_mem_6_cns_csa_n_shi1;
  wire shr_mem_6_cns_csb_n_shi0;
  wire shr_mem_6_cns_csb_n_shi1;
  wire [63:0] shr_mem_6_cns_dinb_shi0;
  wire [63:0] shr_mem_6_cns_dinb_shi1;
  wire [63:0] shr_mem_6_cns_douta_sho0;
  wire [63:0] shr_mem_6_cns_douta_sho1;
  wire shr_mem_6_cns_unc_1;
  wire shr_mem_7_cns_R0;
  wire shr_mem_7_cns_R1;
  wire [7:0] shr_mem_7_cns_addra_shi0;
  wire [7:0] shr_mem_7_cns_addra_shi1;
  wire [7:0] shr_mem_7_cns_addrb_shi0;
  wire [7:0] shr_mem_7_cns_addrb_shi1;
  wire shr_mem_7_cns_csa_n_shi0;
  wire shr_mem_7_cns_csa_n_shi1;
  wire shr_mem_7_cns_csb_n_shi0;
  wire shr_mem_7_cns_csb_n_shi1;
  wire [63:0] shr_mem_7_cns_dinb_shi0;
  wire [63:0] shr_mem_7_cns_dinb_shi1;
  wire [63:0] shr_mem_7_cns_douta_sho0;
  wire [63:0] shr_mem_7_cns_douta_sho1;
  wire shr_mem_7_cns_unc_1;
  wire shr_mem_8_cns_R0;
  wire shr_mem_8_cns_R1;
  wire [7:0] shr_mem_8_cns_addra_shi0;
  wire [7:0] shr_mem_8_cns_addra_shi1;
  wire [7:0] shr_mem_8_cns_addrb_shi0;
  wire [7:0] shr_mem_8_cns_addrb_shi1;
  wire shr_mem_8_cns_csa_n_shi0;
  wire shr_mem_8_cns_csa_n_shi1;
  wire shr_mem_8_cns_csb_n_shi0;
  wire shr_mem_8_cns_csb_n_shi1;
  wire [63:0] shr_mem_8_cns_dinb_shi0;
  wire [63:0] shr_mem_8_cns_dinb_shi1;
  wire [63:0] shr_mem_8_cns_douta_sho0;
  wire [63:0] shr_mem_8_cns_douta_sho1;
  wire shr_mem_8_cns_unc_1;
  wire shr_mem_9_cns_R0;
  wire shr_mem_9_cns_R1;
  wire [7:0] shr_mem_9_cns_addra_shi0;
  wire [7:0] shr_mem_9_cns_addra_shi1;
  wire [7:0] shr_mem_9_cns_addrb_shi0;
  wire [7:0] shr_mem_9_cns_addrb_shi1;
  wire shr_mem_9_cns_csa_n_shi0;
  wire shr_mem_9_cns_csa_n_shi1;
  wire shr_mem_9_cns_csb_n_shi0;
  wire shr_mem_9_cns_csb_n_shi1;
  wire [63:0] shr_mem_9_cns_dinb_shi0;
  wire [63:0] shr_mem_9_cns_dinb_shi1;
  wire [63:0] shr_mem_9_cns_douta_sho0;
  wire [63:0] shr_mem_9_cns_douta_sho1;
  wire shr_mem_9_cns_unc_1;
  wire shr_mem_10_cns_R0;
  wire shr_mem_10_cns_R1;
  wire [7:0] shr_mem_10_cns_addra_shi0;
  wire [7:0] shr_mem_10_cns_addra_shi1;
  wire [7:0] shr_mem_10_cns_addrb_shi0;
  wire [7:0] shr_mem_10_cns_addrb_shi1;
  wire shr_mem_10_cns_csa_n_shi0;
  wire shr_mem_10_cns_csa_n_shi1;
  wire shr_mem_10_cns_csb_n_shi0;
  wire shr_mem_10_cns_csb_n_shi1;
  wire [63:0] shr_mem_10_cns_dinb_shi0;
  wire [63:0] shr_mem_10_cns_dinb_shi1;
  wire [63:0] shr_mem_10_cns_douta_sho0;
  wire [63:0] shr_mem_10_cns_douta_sho1;
  wire shr_mem_10_cns_unc_1;
  wire shr_mem_11_cns_R0;
  wire shr_mem_11_cns_R1;
  wire [7:0] shr_mem_11_cns_addra_shi0;
  wire [7:0] shr_mem_11_cns_addra_shi1;
  wire [7:0] shr_mem_11_cns_addrb_shi0;
  wire [7:0] shr_mem_11_cns_addrb_shi1;
  wire shr_mem_11_cns_csa_n_shi0;
  wire shr_mem_11_cns_csa_n_shi1;
  wire shr_mem_11_cns_csb_n_shi0;
  wire shr_mem_11_cns_csb_n_shi1;
  wire [63:0] shr_mem_11_cns_dinb_shi0;
  wire [63:0] shr_mem_11_cns_dinb_shi1;
  wire [63:0] shr_mem_11_cns_douta_sho0;
  wire [63:0] shr_mem_11_cns_douta_sho1;
  wire shr_mem_11_cns_unc_1;
  wire shr_mem_12_cns_R0;
  wire shr_mem_12_cns_R1;
  wire [7:0] shr_mem_12_cns_addra_shi0;
  wire [7:0] shr_mem_12_cns_addra_shi1;
  wire [7:0] shr_mem_12_cns_addrb_shi0;
  wire [7:0] shr_mem_12_cns_addrb_shi1;
  wire shr_mem_12_cns_csa_n_shi0;
  wire shr_mem_12_cns_csa_n_shi1;
  wire shr_mem_12_cns_csb_n_shi0;
  wire shr_mem_12_cns_csb_n_shi1;
  wire [63:0] shr_mem_12_cns_dinb_shi0;
  wire [63:0] shr_mem_12_cns_dinb_shi1;
  wire [63:0] shr_mem_12_cns_douta_sho0;
  wire [63:0] shr_mem_12_cns_douta_sho1;
  wire shr_mem_12_cns_unc_1;
  wire shr_mem_13_cns_R0;
  wire shr_mem_13_cns_R1;
  wire [7:0] shr_mem_13_cns_addra_shi0;
  wire [7:0] shr_mem_13_cns_addra_shi1;
  wire [7:0] shr_mem_13_cns_addrb_shi0;
  wire [7:0] shr_mem_13_cns_addrb_shi1;
  wire shr_mem_13_cns_csa_n_shi0;
  wire shr_mem_13_cns_csa_n_shi1;
  wire shr_mem_13_cns_csb_n_shi0;
  wire shr_mem_13_cns_csb_n_shi1;
  wire [63:0] shr_mem_13_cns_dinb_shi0;
  wire [63:0] shr_mem_13_cns_dinb_shi1;
  wire [63:0] shr_mem_13_cns_douta_sho0;
  wire [63:0] shr_mem_13_cns_douta_sho1;
  wire shr_mem_13_cns_unc_1;
  wire shr_mem_14_cns_R0;
  wire shr_mem_14_cns_R1;
  wire [7:0] shr_mem_14_cns_addra_shi0;
  wire [7:0] shr_mem_14_cns_addra_shi1;
  wire [7:0] shr_mem_14_cns_addrb_shi0;
  wire [7:0] shr_mem_14_cns_addrb_shi1;
  wire shr_mem_14_cns_csa_n_shi0;
  wire shr_mem_14_cns_csa_n_shi1;
  wire shr_mem_14_cns_csb_n_shi0;
  wire shr_mem_14_cns_csb_n_shi1;
  wire [63:0] shr_mem_14_cns_dinb_shi0;
  wire [63:0] shr_mem_14_cns_dinb_shi1;
  wire [63:0] shr_mem_14_cns_douta_sho0;
  wire [63:0] shr_mem_14_cns_douta_sho1;
  wire shr_mem_14_cns_unc_1;
  wire shr_mem_15_cns_R0;
  wire shr_mem_15_cns_R1;
  wire [7:0] shr_mem_15_cns_addra_shi0;
  wire [7:0] shr_mem_15_cns_addra_shi1;
  wire [7:0] shr_mem_15_cns_addrb_shi0;
  wire [7:0] shr_mem_15_cns_addrb_shi1;
  wire shr_mem_15_cns_csa_n_shi0;
  wire shr_mem_15_cns_csa_n_shi1;
  wire shr_mem_15_cns_csb_n_shi0;
  wire shr_mem_15_cns_csb_n_shi1;
  wire [63:0] shr_mem_15_cns_dinb_shi0;
  wire [63:0] shr_mem_15_cns_dinb_shi1;
  wire [63:0] shr_mem_15_cns_douta_sho0;
  wire [63:0] shr_mem_15_cns_douta_sho1;
  wire shr_mem_15_cns_unc_1;
  wire shr_mem_0_cns_S1_iff;
  wire shr_mem_0_cns_S0_iff;
  wire shr_mem_1_cns_S1_iff;
  wire din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_1_cns_S0_iff;
  wire shr_mem_2_cns_S1_iff;
  wire din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_2_cns_S0_iff;
  wire shr_mem_3_cns_S1_iff;
  wire din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_3_cns_S0_iff;
  wire shr_mem_4_cns_S1_iff;
  wire din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_4_cns_S0_iff;
  wire shr_mem_5_cns_S1_iff;
  wire din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_5_cns_S0_iff;
  wire shr_mem_6_cns_S1_iff;
  wire din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_6_cns_S0_iff;
  wire shr_mem_7_cns_S1_iff;
  wire din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_7_cns_S0_iff;
  wire shr_mem_8_cns_S1_iff;
  wire din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_8_cns_S0_iff;
  wire shr_mem_9_cns_S1_iff;
  wire din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_9_cns_S0_iff;
  wire shr_mem_10_cns_S1_iff;
  wire din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_10_cns_S0_iff;
  wire shr_mem_11_cns_S1_iff;
  wire din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_11_cns_S0_iff;
  wire shr_mem_12_cns_S1_iff;
  wire din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_12_cns_S0_iff;
  wire shr_mem_13_cns_S1_iff;
  wire din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_13_cns_S0_iff;
  wire shr_mem_14_cns_S1_iff;
  wire din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_14_cns_S0_iff;
  wire shr_mem_15_cns_S1_iff;
  wire din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff;
  wire dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff;
  wire shr_mem_15_cns_S0_iff;
  wire shr_mem_0_cns_S0_dmo;
  wire shr_mem_0_cns_S1_dmo;
  wire shr_mem_1_cns_S0_dmo;
  wire shr_mem_1_cns_S1_dmo;
  wire shr_mem_2_cns_S0_dmo;
  wire shr_mem_2_cns_S1_dmo;
  wire shr_mem_3_cns_S0_dmo;
  wire shr_mem_3_cns_S1_dmo;
  wire shr_mem_4_cns_S0_dmo;
  wire shr_mem_4_cns_S1_dmo;
  wire shr_mem_5_cns_S0_dmo;
  wire shr_mem_5_cns_S1_dmo;
  wire shr_mem_6_cns_S0_dmo;
  wire shr_mem_6_cns_S1_dmo;
  wire shr_mem_7_cns_S0_dmo;
  wire shr_mem_7_cns_S1_dmo;
  wire shr_mem_8_cns_S0_dmo;
  wire shr_mem_8_cns_S1_dmo;
  wire shr_mem_9_cns_S0_dmo;
  wire shr_mem_9_cns_S1_dmo;
  wire shr_mem_10_cns_S0_dmo;
  wire shr_mem_10_cns_S1_dmo;
  wire shr_mem_11_cns_S0_dmo;
  wire shr_mem_11_cns_S1_dmo;
  wire shr_mem_12_cns_S0_dmo;
  wire shr_mem_12_cns_S1_dmo;
  wire shr_mem_13_cns_S0_dmo;
  wire shr_mem_13_cns_S1_dmo;
  wire shr_mem_14_cns_S0_dmo;
  wire shr_mem_14_cns_S1_dmo;
  wire shr_mem_15_cns_S0_dmo;
  wire shr_mem_15_cns_S1_dmo;


  // Interconnect Declarations for Component Instantiations 
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_0_cns_comp (
      .addra(shr_mem_0_cns_addra_shi0),
      .addrb(shr_mem_0_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_0_cns_csa_n_shi0),
      .csb_n(shr_mem_0_cns_csb_n_shi0),
      .dinb(shr_mem_0_cns_dinb_shi0),
      .douta(shr_mem_0_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_0_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_0_cns_comp_1 (
      .addra(shr_mem_0_cns_addra_shi1),
      .addrb(shr_mem_0_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_0_cns_csa_n_shi1),
      .csb_n(shr_mem_0_cns_csb_n_shi1),
      .dinb(shr_mem_0_cns_dinb_shi1),
      .douta(shr_mem_0_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_0_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_1_cns_comp (
      .addra(shr_mem_1_cns_addra_shi0),
      .addrb(shr_mem_1_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_1_cns_csa_n_shi0),
      .csb_n(shr_mem_1_cns_csb_n_shi0),
      .dinb(shr_mem_1_cns_dinb_shi0),
      .douta(shr_mem_1_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_1_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_1_cns_comp_1 (
      .addra(shr_mem_1_cns_addra_shi1),
      .addrb(shr_mem_1_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_1_cns_csa_n_shi1),
      .csb_n(shr_mem_1_cns_csb_n_shi1),
      .dinb(shr_mem_1_cns_dinb_shi1),
      .douta(shr_mem_1_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_1_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_2_cns_comp (
      .addra(shr_mem_2_cns_addra_shi0),
      .addrb(shr_mem_2_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_2_cns_csa_n_shi0),
      .csb_n(shr_mem_2_cns_csb_n_shi0),
      .dinb(shr_mem_2_cns_dinb_shi0),
      .douta(shr_mem_2_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_2_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_2_cns_comp_1 (
      .addra(shr_mem_2_cns_addra_shi1),
      .addrb(shr_mem_2_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_2_cns_csa_n_shi1),
      .csb_n(shr_mem_2_cns_csb_n_shi1),
      .dinb(shr_mem_2_cns_dinb_shi1),
      .douta(shr_mem_2_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_2_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_3_cns_comp (
      .addra(shr_mem_3_cns_addra_shi0),
      .addrb(shr_mem_3_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_3_cns_csa_n_shi0),
      .csb_n(shr_mem_3_cns_csb_n_shi0),
      .dinb(shr_mem_3_cns_dinb_shi0),
      .douta(shr_mem_3_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_3_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_3_cns_comp_1 (
      .addra(shr_mem_3_cns_addra_shi1),
      .addrb(shr_mem_3_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_3_cns_csa_n_shi1),
      .csb_n(shr_mem_3_cns_csb_n_shi1),
      .dinb(shr_mem_3_cns_dinb_shi1),
      .douta(shr_mem_3_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_3_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_4_cns_comp (
      .addra(shr_mem_4_cns_addra_shi0),
      .addrb(shr_mem_4_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_4_cns_csa_n_shi0),
      .csb_n(shr_mem_4_cns_csb_n_shi0),
      .dinb(shr_mem_4_cns_dinb_shi0),
      .douta(shr_mem_4_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_4_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_4_cns_comp_1 (
      .addra(shr_mem_4_cns_addra_shi1),
      .addrb(shr_mem_4_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_4_cns_csa_n_shi1),
      .csb_n(shr_mem_4_cns_csb_n_shi1),
      .dinb(shr_mem_4_cns_dinb_shi1),
      .douta(shr_mem_4_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_4_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_5_cns_comp (
      .addra(shr_mem_5_cns_addra_shi0),
      .addrb(shr_mem_5_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_5_cns_csa_n_shi0),
      .csb_n(shr_mem_5_cns_csb_n_shi0),
      .dinb(shr_mem_5_cns_dinb_shi0),
      .douta(shr_mem_5_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_5_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_5_cns_comp_1 (
      .addra(shr_mem_5_cns_addra_shi1),
      .addrb(shr_mem_5_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_5_cns_csa_n_shi1),
      .csb_n(shr_mem_5_cns_csb_n_shi1),
      .dinb(shr_mem_5_cns_dinb_shi1),
      .douta(shr_mem_5_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_5_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_6_cns_comp (
      .addra(shr_mem_6_cns_addra_shi0),
      .addrb(shr_mem_6_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_6_cns_csa_n_shi0),
      .csb_n(shr_mem_6_cns_csb_n_shi0),
      .dinb(shr_mem_6_cns_dinb_shi0),
      .douta(shr_mem_6_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_6_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_6_cns_comp_1 (
      .addra(shr_mem_6_cns_addra_shi1),
      .addrb(shr_mem_6_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_6_cns_csa_n_shi1),
      .csb_n(shr_mem_6_cns_csb_n_shi1),
      .dinb(shr_mem_6_cns_dinb_shi1),
      .douta(shr_mem_6_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_6_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_7_cns_comp (
      .addra(shr_mem_7_cns_addra_shi0),
      .addrb(shr_mem_7_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_7_cns_csa_n_shi0),
      .csb_n(shr_mem_7_cns_csb_n_shi0),
      .dinb(shr_mem_7_cns_dinb_shi0),
      .douta(shr_mem_7_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_7_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_7_cns_comp_1 (
      .addra(shr_mem_7_cns_addra_shi1),
      .addrb(shr_mem_7_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_7_cns_csa_n_shi1),
      .csb_n(shr_mem_7_cns_csb_n_shi1),
      .dinb(shr_mem_7_cns_dinb_shi1),
      .douta(shr_mem_7_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_7_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_8_cns_comp (
      .addra(shr_mem_8_cns_addra_shi0),
      .addrb(shr_mem_8_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_8_cns_csa_n_shi0),
      .csb_n(shr_mem_8_cns_csb_n_shi0),
      .dinb(shr_mem_8_cns_dinb_shi0),
      .douta(shr_mem_8_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_8_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_8_cns_comp_1 (
      .addra(shr_mem_8_cns_addra_shi1),
      .addrb(shr_mem_8_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_8_cns_csa_n_shi1),
      .csb_n(shr_mem_8_cns_csb_n_shi1),
      .dinb(shr_mem_8_cns_dinb_shi1),
      .douta(shr_mem_8_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_8_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_9_cns_comp (
      .addra(shr_mem_9_cns_addra_shi0),
      .addrb(shr_mem_9_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_9_cns_csa_n_shi0),
      .csb_n(shr_mem_9_cns_csb_n_shi0),
      .dinb(shr_mem_9_cns_dinb_shi0),
      .douta(shr_mem_9_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_9_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_9_cns_comp_1 (
      .addra(shr_mem_9_cns_addra_shi1),
      .addrb(shr_mem_9_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_9_cns_csa_n_shi1),
      .csb_n(shr_mem_9_cns_csb_n_shi1),
      .dinb(shr_mem_9_cns_dinb_shi1),
      .douta(shr_mem_9_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_9_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_10_cns_comp (
      .addra(shr_mem_10_cns_addra_shi0),
      .addrb(shr_mem_10_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_10_cns_csa_n_shi0),
      .csb_n(shr_mem_10_cns_csb_n_shi0),
      .dinb(shr_mem_10_cns_dinb_shi0),
      .douta(shr_mem_10_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_10_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_10_cns_comp_1 (
      .addra(shr_mem_10_cns_addra_shi1),
      .addrb(shr_mem_10_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_10_cns_csa_n_shi1),
      .csb_n(shr_mem_10_cns_csb_n_shi1),
      .dinb(shr_mem_10_cns_dinb_shi1),
      .douta(shr_mem_10_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_10_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_11_cns_comp (
      .addra(shr_mem_11_cns_addra_shi0),
      .addrb(shr_mem_11_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_11_cns_csa_n_shi0),
      .csb_n(shr_mem_11_cns_csb_n_shi0),
      .dinb(shr_mem_11_cns_dinb_shi0),
      .douta(shr_mem_11_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_11_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_11_cns_comp_1 (
      .addra(shr_mem_11_cns_addra_shi1),
      .addrb(shr_mem_11_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_11_cns_csa_n_shi1),
      .csb_n(shr_mem_11_cns_csb_n_shi1),
      .dinb(shr_mem_11_cns_dinb_shi1),
      .douta(shr_mem_11_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_11_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_12_cns_comp (
      .addra(shr_mem_12_cns_addra_shi0),
      .addrb(shr_mem_12_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_12_cns_csa_n_shi0),
      .csb_n(shr_mem_12_cns_csb_n_shi0),
      .dinb(shr_mem_12_cns_dinb_shi0),
      .douta(shr_mem_12_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_12_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_12_cns_comp_1 (
      .addra(shr_mem_12_cns_addra_shi1),
      .addrb(shr_mem_12_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_12_cns_csa_n_shi1),
      .csb_n(shr_mem_12_cns_csb_n_shi1),
      .dinb(shr_mem_12_cns_dinb_shi1),
      .douta(shr_mem_12_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_12_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_13_cns_comp (
      .addra(shr_mem_13_cns_addra_shi0),
      .addrb(shr_mem_13_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_13_cns_csa_n_shi0),
      .csb_n(shr_mem_13_cns_csb_n_shi0),
      .dinb(shr_mem_13_cns_dinb_shi0),
      .douta(shr_mem_13_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_13_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_13_cns_comp_1 (
      .addra(shr_mem_13_cns_addra_shi1),
      .addrb(shr_mem_13_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_13_cns_csa_n_shi1),
      .csb_n(shr_mem_13_cns_csb_n_shi1),
      .dinb(shr_mem_13_cns_dinb_shi1),
      .douta(shr_mem_13_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_13_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_14_cns_comp (
      .addra(shr_mem_14_cns_addra_shi0),
      .addrb(shr_mem_14_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_14_cns_csa_n_shi0),
      .csb_n(shr_mem_14_cns_csb_n_shi0),
      .dinb(shr_mem_14_cns_dinb_shi0),
      .douta(shr_mem_14_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_14_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_14_cns_comp_1 (
      .addra(shr_mem_14_cns_addra_shi1),
      .addrb(shr_mem_14_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_14_cns_csa_n_shi1),
      .csb_n(shr_mem_14_cns_csb_n_shi1),
      .dinb(shr_mem_14_cns_dinb_shi1),
      .douta(shr_mem_14_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_14_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_15_cns_comp (
      .addra(shr_mem_15_cns_addra_shi0),
      .addrb(shr_mem_15_cns_addrb_shi0),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_15_cns_csa_n_shi0),
      .csb_n(shr_mem_15_cns_csb_n_shi0),
      .dinb(shr_mem_15_cns_dinb_shi0),
      .douta(shr_mem_15_cns_douta_sho0),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_15_cns_unc_1)
    );
  cat_ram2p_half #(.filename(-1073740000),
  .MEMORY_ACC_WIDTH(-1073740000)) shr_mem_15_cns_comp_1 (
      .addra(shr_mem_15_cns_addra_shi1),
      .addrb(shr_mem_15_cns_addrb_shi1),
      .clamp_mem(clamp_mem),
      .clk(clk),
      .csa_n(shr_mem_15_cns_csa_n_shi1),
      .csb_n(shr_mem_15_cns_csb_n_shi1),
      .dinb(shr_mem_15_cns_dinb_shi1),
      .douta(shr_mem_15_cns_douta_sho1),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .sin(1'b0),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n),
      .sout(shr_mem_15_cns_unc_1)
    );
  WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_1 WRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(din_rsc_z),
      .din_rsc_vz(din_rsc_vz),
      .din_rsc_lz(din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_0_rsc_csa_n(dout_0_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_csb_n(dout_0_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_addra(dout_0_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_addrb(dout_0_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_dinb(dout_0_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_douta(dout_0_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_req_vz(dout_0_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_rls_lz(dout_0_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_1_rsc_csa_n(dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_csb_n(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_addra(dout_1_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_addrb(dout_1_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_dinb(dout_1_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_douta(dout_1_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_req_vz(dout_1_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_rls_lz(dout_1_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_2_rsc_csa_n(dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_csb_n(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_addra(dout_2_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_addrb(dout_2_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_dinb(dout_2_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_douta(dout_2_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_req_vz(dout_2_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_rls_lz(dout_2_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_3_rsc_csa_n(dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_csb_n(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_addra(dout_3_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_addrb(dout_3_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_dinb(dout_3_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_douta(dout_3_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_req_vz(dout_3_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_rls_lz(dout_3_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_4_rsc_csa_n(dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_csb_n(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_addra(dout_4_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_addrb(dout_4_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_dinb(dout_4_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_douta(dout_4_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_req_vz(dout_4_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_rls_lz(dout_4_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_5_rsc_csa_n(dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_csb_n(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_addra(dout_5_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_addrb(dout_5_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_dinb(dout_5_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_douta(dout_5_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_req_vz(dout_5_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_rls_lz(dout_5_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_6_rsc_csa_n(dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_csb_n(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_addra(dout_6_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_addrb(dout_6_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_dinb(dout_6_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_douta(dout_6_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_req_vz(dout_6_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_rls_lz(dout_6_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_7_rsc_csa_n(dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_csb_n(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_addra(dout_7_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_addrb(dout_7_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_dinb(dout_7_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_douta(dout_7_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_req_vz(dout_7_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_rls_lz(dout_7_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_8_rsc_csa_n(dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_csb_n(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_addra(dout_8_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_addrb(dout_8_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_dinb(dout_8_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_douta(dout_8_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_req_vz(dout_8_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_rls_lz(dout_8_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_9_rsc_csa_n(dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_csb_n(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_addra(dout_9_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_addrb(dout_9_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_dinb(dout_9_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_douta(dout_9_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_req_vz(dout_9_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_rls_lz(dout_9_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_10_rsc_csa_n(dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_csb_n(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_addra(dout_10_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_addrb(dout_10_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_dinb(dout_10_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_douta(dout_10_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_req_vz(dout_10_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_rls_lz(dout_10_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_11_rsc_csa_n(dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_csb_n(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_addra(dout_11_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_addrb(dout_11_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_dinb(dout_11_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_douta(dout_11_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_req_vz(dout_11_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_rls_lz(dout_11_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_12_rsc_csa_n(dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_csb_n(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_addra(dout_12_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_addrb(dout_12_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_dinb(dout_12_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_douta(dout_12_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_req_vz(dout_12_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_rls_lz(dout_12_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_13_rsc_csa_n(dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_csb_n(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_addra(dout_13_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_addrb(dout_13_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_dinb(dout_13_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_douta(dout_13_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_req_vz(dout_13_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_rls_lz(dout_13_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_14_rsc_csa_n(dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_csb_n(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_addra(dout_14_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_addrb(dout_14_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_dinb(dout_14_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_douta(dout_14_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_req_vz(dout_14_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_rls_lz(dout_14_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_15_rsc_csa_n(dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_csb_n(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_addra(dout_15_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_addrb(dout_15_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_dinb(dout_15_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_douta(dout_15_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_req_vz(dout_15_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_rls_lz(dout_15_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud)
    );
  READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_1 READ_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst (
      .clk(clk),
      .rst(rst),
      .din_0_rsc_csa_n(din_0_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_csb_n(din_0_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_addra(din_0_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_addrb(din_0_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_dinb(din_0_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_douta(din_0_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_req_vz(din_0_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_rls_lz(din_0_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_1_rsc_csa_n(din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_csb_n(din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_addra(din_1_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_addrb(din_1_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_dinb(din_1_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_douta(din_1_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_req_vz(din_1_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_rls_lz(din_1_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_2_rsc_csa_n(din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_csb_n(din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_addra(din_2_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_addrb(din_2_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_dinb(din_2_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_douta(din_2_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_req_vz(din_2_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_rls_lz(din_2_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_3_rsc_csa_n(din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_csb_n(din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_addra(din_3_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_addrb(din_3_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_dinb(din_3_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_douta(din_3_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_req_vz(din_3_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_rls_lz(din_3_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_4_rsc_csa_n(din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_csb_n(din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_addra(din_4_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_addrb(din_4_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_dinb(din_4_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_douta(din_4_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_req_vz(din_4_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_rls_lz(din_4_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_5_rsc_csa_n(din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_csb_n(din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_addra(din_5_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_addrb(din_5_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_dinb(din_5_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_douta(din_5_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_req_vz(din_5_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_rls_lz(din_5_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_6_rsc_csa_n(din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_csb_n(din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_addra(din_6_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_addrb(din_6_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_dinb(din_6_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_douta(din_6_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_req_vz(din_6_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_rls_lz(din_6_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_7_rsc_csa_n(din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_csb_n(din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_addra(din_7_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_addrb(din_7_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_dinb(din_7_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_douta(din_7_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_req_vz(din_7_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_rls_lz(din_7_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_8_rsc_csa_n(din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_csb_n(din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_addra(din_8_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_addrb(din_8_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_dinb(din_8_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_douta(din_8_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_req_vz(din_8_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_rls_lz(din_8_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_9_rsc_csa_n(din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_csb_n(din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_addra(din_9_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_addrb(din_9_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_dinb(din_9_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_douta(din_9_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_req_vz(din_9_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_rls_lz(din_9_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_10_rsc_csa_n(din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_csb_n(din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_addra(din_10_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_addrb(din_10_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_dinb(din_10_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_douta(din_10_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_req_vz(din_10_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_rls_lz(din_10_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_11_rsc_csa_n(din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_csb_n(din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_addra(din_11_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_addrb(din_11_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_dinb(din_11_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_douta(din_11_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_req_vz(din_11_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_rls_lz(din_11_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_12_rsc_csa_n(din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_csb_n(din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_addra(din_12_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_addrb(din_12_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_dinb(din_12_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_douta(din_12_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_req_vz(din_12_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_rls_lz(din_12_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_13_rsc_csa_n(din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_csb_n(din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_addra(din_13_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_addrb(din_13_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_dinb(din_13_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_douta(din_13_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_req_vz(din_13_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_rls_lz(din_13_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_14_rsc_csa_n(din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_csb_n(din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_addra(din_14_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_addrb(din_14_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_dinb(din_14_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_douta(din_14_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_req_vz(din_14_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_rls_lz(din_14_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_15_rsc_csa_n(din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_csb_n(din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_addra(din_15_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_addrb(din_15_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_dinb(din_15_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_douta(din_15_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_req_vz(din_15_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_rls_lz(din_15_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_rsc_z(dout_rsc_z_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_rsc_vz(dout_rsc_vz),
      .dout_rsc_lz(dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud)
    );
  unreg_hier_31 unreg (
      .in_0(shr_mem_0_cns_S0_iff),
      .out_0(shr_mem_0_cns_R0)
    );
  unreg_hier_31 unreg_1 (
      .in_0(shr_mem_0_cns_S1_iff),
      .out_0(shr_mem_0_cns_R1)
    );
  unreg_hier_31 unreg_2 (
      .in_0(shr_mem_1_cns_S0_iff),
      .out_0(shr_mem_1_cns_R0)
    );
  unreg_hier_31 unreg_3 (
      .in_0(shr_mem_1_cns_S1_iff),
      .out_0(shr_mem_1_cns_R1)
    );
  unreg_hier_31 unreg_4 (
      .in_0(shr_mem_2_cns_S0_iff),
      .out_0(shr_mem_2_cns_R0)
    );
  unreg_hier_31 unreg_5 (
      .in_0(shr_mem_2_cns_S1_iff),
      .out_0(shr_mem_2_cns_R1)
    );
  unreg_hier_31 unreg_6 (
      .in_0(shr_mem_3_cns_S0_iff),
      .out_0(shr_mem_3_cns_R0)
    );
  unreg_hier_31 unreg_7 (
      .in_0(shr_mem_3_cns_S1_iff),
      .out_0(shr_mem_3_cns_R1)
    );
  unreg_hier_31 unreg_8 (
      .in_0(shr_mem_4_cns_S0_iff),
      .out_0(shr_mem_4_cns_R0)
    );
  unreg_hier_31 unreg_9 (
      .in_0(shr_mem_4_cns_S1_iff),
      .out_0(shr_mem_4_cns_R1)
    );
  unreg_hier_31 unreg_10 (
      .in_0(shr_mem_5_cns_S0_iff),
      .out_0(shr_mem_5_cns_R0)
    );
  unreg_hier_31 unreg_11 (
      .in_0(shr_mem_5_cns_S1_iff),
      .out_0(shr_mem_5_cns_R1)
    );
  unreg_hier_31 unreg_12 (
      .in_0(shr_mem_6_cns_S0_iff),
      .out_0(shr_mem_6_cns_R0)
    );
  unreg_hier_31 unreg_13 (
      .in_0(shr_mem_6_cns_S1_iff),
      .out_0(shr_mem_6_cns_R1)
    );
  unreg_hier_31 unreg_14 (
      .in_0(shr_mem_7_cns_S0_iff),
      .out_0(shr_mem_7_cns_R0)
    );
  unreg_hier_31 unreg_15 (
      .in_0(shr_mem_7_cns_S1_iff),
      .out_0(shr_mem_7_cns_R1)
    );
  unreg_hier_31 unreg_16 (
      .in_0(shr_mem_8_cns_S0_iff),
      .out_0(shr_mem_8_cns_R0)
    );
  unreg_hier_31 unreg_17 (
      .in_0(shr_mem_8_cns_S1_iff),
      .out_0(shr_mem_8_cns_R1)
    );
  unreg_hier_31 unreg_18 (
      .in_0(shr_mem_9_cns_S0_iff),
      .out_0(shr_mem_9_cns_R0)
    );
  unreg_hier_31 unreg_19 (
      .in_0(shr_mem_9_cns_S1_iff),
      .out_0(shr_mem_9_cns_R1)
    );
  unreg_hier_31 unreg_20 (
      .in_0(shr_mem_10_cns_S0_iff),
      .out_0(shr_mem_10_cns_R0)
    );
  unreg_hier_31 unreg_21 (
      .in_0(shr_mem_10_cns_S1_iff),
      .out_0(shr_mem_10_cns_R1)
    );
  unreg_hier_31 unreg_22 (
      .in_0(shr_mem_11_cns_S0_iff),
      .out_0(shr_mem_11_cns_R0)
    );
  unreg_hier_31 unreg_23 (
      .in_0(shr_mem_11_cns_S1_iff),
      .out_0(shr_mem_11_cns_R1)
    );
  unreg_hier_31 unreg_24 (
      .in_0(shr_mem_12_cns_S0_iff),
      .out_0(shr_mem_12_cns_R0)
    );
  unreg_hier_31 unreg_25 (
      .in_0(shr_mem_12_cns_S1_iff),
      .out_0(shr_mem_12_cns_R1)
    );
  unreg_hier_31 unreg_26 (
      .in_0(shr_mem_13_cns_S0_iff),
      .out_0(shr_mem_13_cns_R0)
    );
  unreg_hier_31 unreg_27 (
      .in_0(shr_mem_13_cns_S1_iff),
      .out_0(shr_mem_13_cns_R1)
    );
  unreg_hier_31 unreg_28 (
      .in_0(shr_mem_14_cns_S0_iff),
      .out_0(shr_mem_14_cns_R0)
    );
  unreg_hier_31 unreg_29 (
      .in_0(shr_mem_14_cns_S1_iff),
      .out_0(shr_mem_14_cns_R1)
    );
  unreg_hier_31 unreg_30 (
      .in_0(shr_mem_15_cns_S0_iff),
      .out_0(shr_mem_15_cns_R0)
    );
  unreg_hier_31 unreg_31 (
      .in_0(shr_mem_15_cns_S1_iff),
      .out_0(shr_mem_15_cns_R1)
    );
  double_buffeYeetf_0_cns_bctl double_buffeYeetf_0_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(1'b0),
      .dout_0_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_0_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_0_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_0_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_0_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_0_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_0_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_0_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_0_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(1'b0),
      .din_0_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_0_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_0_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_0_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_0_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_0_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_0_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_0_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz),
      .din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_0_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_0_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_0_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_0_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_1_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_1_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_2_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_2_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_3_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_3_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_4_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_4_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_5_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_5_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_6_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_6_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_7_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_7_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_8_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_8_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_9_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_9_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_10_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_10_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_11_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_11_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_12_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_12_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_13_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_13_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_14_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_14_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .dout_15_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(1'b0),
      .din_15_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(1'b0),
      .dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_0_cns_S0(shr_mem_0_cns_S0_dmo),
      .shr_mem_0_cns_R0(shr_mem_0_cns_R0),
      .shr_mem_0_cns_S1(shr_mem_0_cns_S1_dmo),
      .shr_mem_0_cns_R1(shr_mem_0_cns_R1),
      .shr_mem_0_cns_addra_shi0(shr_mem_0_cns_addra_shi0),
      .shr_mem_0_cns_addra_shi1(shr_mem_0_cns_addra_shi1),
      .shr_mem_0_cns_addrb_shi0(shr_mem_0_cns_addrb_shi0),
      .shr_mem_0_cns_addrb_shi1(shr_mem_0_cns_addrb_shi1),
      .shr_mem_0_cns_csa_n_shi0(shr_mem_0_cns_csa_n_shi0),
      .shr_mem_0_cns_csa_n_shi1(shr_mem_0_cns_csa_n_shi1),
      .shr_mem_0_cns_csb_n_shi0(shr_mem_0_cns_csb_n_shi0),
      .shr_mem_0_cns_csb_n_shi1(shr_mem_0_cns_csb_n_shi1),
      .shr_mem_0_cns_dinb_shi0(shr_mem_0_cns_dinb_shi0),
      .shr_mem_0_cns_dinb_shi1(shr_mem_0_cns_dinb_shi1),
      .shr_mem_0_cns_douta_sho0(shr_mem_0_cns_douta_sho0),
      .shr_mem_0_cns_douta_sho1(shr_mem_0_cns_douta_sho1),
      .shr_mem_0_cns_S1_pff(shr_mem_0_cns_S1_iff),
      .shr_mem_0_cns_S0_pff(shr_mem_0_cns_S0_iff),
      .din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff)
    );
  double_buffeYeetf_1_cns_bctl double_buffeYeetf_1_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_1_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_1_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_1_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_1_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_1_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_1_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_1_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_1_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_1_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_1_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_1_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_1_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_1_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_1_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_1_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_1_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_1_cns_S0(shr_mem_1_cns_S0_dmo),
      .shr_mem_1_cns_R0(shr_mem_1_cns_R0),
      .shr_mem_1_cns_S1(shr_mem_1_cns_S1_dmo),
      .shr_mem_1_cns_R1(shr_mem_1_cns_R1),
      .shr_mem_1_cns_addra_shi0(shr_mem_1_cns_addra_shi0),
      .shr_mem_1_cns_addra_shi1(shr_mem_1_cns_addra_shi1),
      .shr_mem_1_cns_addrb_shi0(shr_mem_1_cns_addrb_shi0),
      .shr_mem_1_cns_addrb_shi1(shr_mem_1_cns_addrb_shi1),
      .shr_mem_1_cns_csa_n_shi0(shr_mem_1_cns_csa_n_shi0),
      .shr_mem_1_cns_csa_n_shi1(shr_mem_1_cns_csa_n_shi1),
      .shr_mem_1_cns_csb_n_shi0(shr_mem_1_cns_csb_n_shi0),
      .shr_mem_1_cns_csb_n_shi1(shr_mem_1_cns_csb_n_shi1),
      .shr_mem_1_cns_dinb_shi0(shr_mem_1_cns_dinb_shi0),
      .shr_mem_1_cns_dinb_shi1(shr_mem_1_cns_dinb_shi1),
      .shr_mem_1_cns_douta_sho0(shr_mem_1_cns_douta_sho0),
      .shr_mem_1_cns_douta_sho1(shr_mem_1_cns_douta_sho1),
      .shr_mem_1_cns_S1_pff(shr_mem_1_cns_S1_iff),
      .din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_1_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_1_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_1_cns_S0_pff(shr_mem_1_cns_S0_iff)
    );
  double_buffeYeetf_2_cns_bctl double_buffeYeetf_2_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_2_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_2_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_2_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_2_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_2_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_2_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_2_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_2_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_2_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_2_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_2_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_2_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_2_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_2_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_2_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_2_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_2_cns_S0(shr_mem_2_cns_S0_dmo),
      .shr_mem_2_cns_R0(shr_mem_2_cns_R0),
      .shr_mem_2_cns_S1(shr_mem_2_cns_S1_dmo),
      .shr_mem_2_cns_R1(shr_mem_2_cns_R1),
      .shr_mem_2_cns_addra_shi0(shr_mem_2_cns_addra_shi0),
      .shr_mem_2_cns_addra_shi1(shr_mem_2_cns_addra_shi1),
      .shr_mem_2_cns_addrb_shi0(shr_mem_2_cns_addrb_shi0),
      .shr_mem_2_cns_addrb_shi1(shr_mem_2_cns_addrb_shi1),
      .shr_mem_2_cns_csa_n_shi0(shr_mem_2_cns_csa_n_shi0),
      .shr_mem_2_cns_csa_n_shi1(shr_mem_2_cns_csa_n_shi1),
      .shr_mem_2_cns_csb_n_shi0(shr_mem_2_cns_csb_n_shi0),
      .shr_mem_2_cns_csb_n_shi1(shr_mem_2_cns_csb_n_shi1),
      .shr_mem_2_cns_dinb_shi0(shr_mem_2_cns_dinb_shi0),
      .shr_mem_2_cns_dinb_shi1(shr_mem_2_cns_dinb_shi1),
      .shr_mem_2_cns_douta_sho0(shr_mem_2_cns_douta_sho0),
      .shr_mem_2_cns_douta_sho1(shr_mem_2_cns_douta_sho1),
      .shr_mem_2_cns_S1_pff(shr_mem_2_cns_S1_iff),
      .din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_2_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_2_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_2_cns_S0_pff(shr_mem_2_cns_S0_iff)
    );
  double_buffeYeetf_3_cns_bctl double_buffeYeetf_3_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_3_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_3_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_3_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_3_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_3_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_3_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_3_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_3_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_3_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_3_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_3_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_3_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_3_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_3_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_3_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_3_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_3_cns_S0(shr_mem_3_cns_S0_dmo),
      .shr_mem_3_cns_R0(shr_mem_3_cns_R0),
      .shr_mem_3_cns_S1(shr_mem_3_cns_S1_dmo),
      .shr_mem_3_cns_R1(shr_mem_3_cns_R1),
      .shr_mem_3_cns_addra_shi0(shr_mem_3_cns_addra_shi0),
      .shr_mem_3_cns_addra_shi1(shr_mem_3_cns_addra_shi1),
      .shr_mem_3_cns_addrb_shi0(shr_mem_3_cns_addrb_shi0),
      .shr_mem_3_cns_addrb_shi1(shr_mem_3_cns_addrb_shi1),
      .shr_mem_3_cns_csa_n_shi0(shr_mem_3_cns_csa_n_shi0),
      .shr_mem_3_cns_csa_n_shi1(shr_mem_3_cns_csa_n_shi1),
      .shr_mem_3_cns_csb_n_shi0(shr_mem_3_cns_csb_n_shi0),
      .shr_mem_3_cns_csb_n_shi1(shr_mem_3_cns_csb_n_shi1),
      .shr_mem_3_cns_dinb_shi0(shr_mem_3_cns_dinb_shi0),
      .shr_mem_3_cns_dinb_shi1(shr_mem_3_cns_dinb_shi1),
      .shr_mem_3_cns_douta_sho0(shr_mem_3_cns_douta_sho0),
      .shr_mem_3_cns_douta_sho1(shr_mem_3_cns_douta_sho1),
      .shr_mem_3_cns_S1_pff(shr_mem_3_cns_S1_iff),
      .din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_3_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_3_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_3_cns_S0_pff(shr_mem_3_cns_S0_iff)
    );
  double_buffeYeetf_4_cns_bctl double_buffeYeetf_4_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_4_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_4_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_4_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_4_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_4_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_4_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_4_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_4_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_4_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_4_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_4_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_4_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_4_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_4_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_4_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_4_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_4_cns_S0(shr_mem_4_cns_S0_dmo),
      .shr_mem_4_cns_R0(shr_mem_4_cns_R0),
      .shr_mem_4_cns_S1(shr_mem_4_cns_S1_dmo),
      .shr_mem_4_cns_R1(shr_mem_4_cns_R1),
      .shr_mem_4_cns_addra_shi0(shr_mem_4_cns_addra_shi0),
      .shr_mem_4_cns_addra_shi1(shr_mem_4_cns_addra_shi1),
      .shr_mem_4_cns_addrb_shi0(shr_mem_4_cns_addrb_shi0),
      .shr_mem_4_cns_addrb_shi1(shr_mem_4_cns_addrb_shi1),
      .shr_mem_4_cns_csa_n_shi0(shr_mem_4_cns_csa_n_shi0),
      .shr_mem_4_cns_csa_n_shi1(shr_mem_4_cns_csa_n_shi1),
      .shr_mem_4_cns_csb_n_shi0(shr_mem_4_cns_csb_n_shi0),
      .shr_mem_4_cns_csb_n_shi1(shr_mem_4_cns_csb_n_shi1),
      .shr_mem_4_cns_dinb_shi0(shr_mem_4_cns_dinb_shi0),
      .shr_mem_4_cns_dinb_shi1(shr_mem_4_cns_dinb_shi1),
      .shr_mem_4_cns_douta_sho0(shr_mem_4_cns_douta_sho0),
      .shr_mem_4_cns_douta_sho1(shr_mem_4_cns_douta_sho1),
      .shr_mem_4_cns_S1_pff(shr_mem_4_cns_S1_iff),
      .din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_4_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_4_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_4_cns_S0_pff(shr_mem_4_cns_S0_iff)
    );
  double_buffeYeetf_5_cns_bctl double_buffeYeetf_5_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_5_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_5_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_5_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_5_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_5_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_5_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_5_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_5_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_5_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_5_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_5_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_5_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_5_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_5_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_5_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_5_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_5_cns_S0(shr_mem_5_cns_S0_dmo),
      .shr_mem_5_cns_R0(shr_mem_5_cns_R0),
      .shr_mem_5_cns_S1(shr_mem_5_cns_S1_dmo),
      .shr_mem_5_cns_R1(shr_mem_5_cns_R1),
      .shr_mem_5_cns_addra_shi0(shr_mem_5_cns_addra_shi0),
      .shr_mem_5_cns_addra_shi1(shr_mem_5_cns_addra_shi1),
      .shr_mem_5_cns_addrb_shi0(shr_mem_5_cns_addrb_shi0),
      .shr_mem_5_cns_addrb_shi1(shr_mem_5_cns_addrb_shi1),
      .shr_mem_5_cns_csa_n_shi0(shr_mem_5_cns_csa_n_shi0),
      .shr_mem_5_cns_csa_n_shi1(shr_mem_5_cns_csa_n_shi1),
      .shr_mem_5_cns_csb_n_shi0(shr_mem_5_cns_csb_n_shi0),
      .shr_mem_5_cns_csb_n_shi1(shr_mem_5_cns_csb_n_shi1),
      .shr_mem_5_cns_dinb_shi0(shr_mem_5_cns_dinb_shi0),
      .shr_mem_5_cns_dinb_shi1(shr_mem_5_cns_dinb_shi1),
      .shr_mem_5_cns_douta_sho0(shr_mem_5_cns_douta_sho0),
      .shr_mem_5_cns_douta_sho1(shr_mem_5_cns_douta_sho1),
      .shr_mem_5_cns_S1_pff(shr_mem_5_cns_S1_iff),
      .din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_5_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_5_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_5_cns_S0_pff(shr_mem_5_cns_S0_iff)
    );
  double_buffeYeetf_6_cns_bctl double_buffeYeetf_6_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_6_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_6_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_6_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_6_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_6_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_6_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_6_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_6_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_6_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_6_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_6_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_6_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_6_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_6_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_6_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_6_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_6_cns_S0(shr_mem_6_cns_S0_dmo),
      .shr_mem_6_cns_R0(shr_mem_6_cns_R0),
      .shr_mem_6_cns_S1(shr_mem_6_cns_S1_dmo),
      .shr_mem_6_cns_R1(shr_mem_6_cns_R1),
      .shr_mem_6_cns_addra_shi0(shr_mem_6_cns_addra_shi0),
      .shr_mem_6_cns_addra_shi1(shr_mem_6_cns_addra_shi1),
      .shr_mem_6_cns_addrb_shi0(shr_mem_6_cns_addrb_shi0),
      .shr_mem_6_cns_addrb_shi1(shr_mem_6_cns_addrb_shi1),
      .shr_mem_6_cns_csa_n_shi0(shr_mem_6_cns_csa_n_shi0),
      .shr_mem_6_cns_csa_n_shi1(shr_mem_6_cns_csa_n_shi1),
      .shr_mem_6_cns_csb_n_shi0(shr_mem_6_cns_csb_n_shi0),
      .shr_mem_6_cns_csb_n_shi1(shr_mem_6_cns_csb_n_shi1),
      .shr_mem_6_cns_dinb_shi0(shr_mem_6_cns_dinb_shi0),
      .shr_mem_6_cns_dinb_shi1(shr_mem_6_cns_dinb_shi1),
      .shr_mem_6_cns_douta_sho0(shr_mem_6_cns_douta_sho0),
      .shr_mem_6_cns_douta_sho1(shr_mem_6_cns_douta_sho1),
      .shr_mem_6_cns_S1_pff(shr_mem_6_cns_S1_iff),
      .din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_6_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_6_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_6_cns_S0_pff(shr_mem_6_cns_S0_iff)
    );
  double_buffeYeetf_7_cns_bctl double_buffeYeetf_7_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_7_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_7_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_7_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_7_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_7_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_7_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_7_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_7_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_7_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_7_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_7_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_7_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_7_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_7_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_7_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_7_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_7_cns_S0(shr_mem_7_cns_S0_dmo),
      .shr_mem_7_cns_R0(shr_mem_7_cns_R0),
      .shr_mem_7_cns_S1(shr_mem_7_cns_S1_dmo),
      .shr_mem_7_cns_R1(shr_mem_7_cns_R1),
      .shr_mem_7_cns_addra_shi0(shr_mem_7_cns_addra_shi0),
      .shr_mem_7_cns_addra_shi1(shr_mem_7_cns_addra_shi1),
      .shr_mem_7_cns_addrb_shi0(shr_mem_7_cns_addrb_shi0),
      .shr_mem_7_cns_addrb_shi1(shr_mem_7_cns_addrb_shi1),
      .shr_mem_7_cns_csa_n_shi0(shr_mem_7_cns_csa_n_shi0),
      .shr_mem_7_cns_csa_n_shi1(shr_mem_7_cns_csa_n_shi1),
      .shr_mem_7_cns_csb_n_shi0(shr_mem_7_cns_csb_n_shi0),
      .shr_mem_7_cns_csb_n_shi1(shr_mem_7_cns_csb_n_shi1),
      .shr_mem_7_cns_dinb_shi0(shr_mem_7_cns_dinb_shi0),
      .shr_mem_7_cns_dinb_shi1(shr_mem_7_cns_dinb_shi1),
      .shr_mem_7_cns_douta_sho0(shr_mem_7_cns_douta_sho0),
      .shr_mem_7_cns_douta_sho1(shr_mem_7_cns_douta_sho1),
      .shr_mem_7_cns_S1_pff(shr_mem_7_cns_S1_iff),
      .din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_7_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_7_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_7_cns_S0_pff(shr_mem_7_cns_S0_iff)
    );
  double_buffeYeetf_8_cns_bctl double_buffeYeetf_8_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_8_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_8_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_8_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_8_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_8_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_8_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_8_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_8_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_8_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_8_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_8_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_8_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_8_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_8_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_8_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_8_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_8_cns_S0(shr_mem_8_cns_S0_dmo),
      .shr_mem_8_cns_R0(shr_mem_8_cns_R0),
      .shr_mem_8_cns_S1(shr_mem_8_cns_S1_dmo),
      .shr_mem_8_cns_R1(shr_mem_8_cns_R1),
      .shr_mem_8_cns_addra_shi0(shr_mem_8_cns_addra_shi0),
      .shr_mem_8_cns_addra_shi1(shr_mem_8_cns_addra_shi1),
      .shr_mem_8_cns_addrb_shi0(shr_mem_8_cns_addrb_shi0),
      .shr_mem_8_cns_addrb_shi1(shr_mem_8_cns_addrb_shi1),
      .shr_mem_8_cns_csa_n_shi0(shr_mem_8_cns_csa_n_shi0),
      .shr_mem_8_cns_csa_n_shi1(shr_mem_8_cns_csa_n_shi1),
      .shr_mem_8_cns_csb_n_shi0(shr_mem_8_cns_csb_n_shi0),
      .shr_mem_8_cns_csb_n_shi1(shr_mem_8_cns_csb_n_shi1),
      .shr_mem_8_cns_dinb_shi0(shr_mem_8_cns_dinb_shi0),
      .shr_mem_8_cns_dinb_shi1(shr_mem_8_cns_dinb_shi1),
      .shr_mem_8_cns_douta_sho0(shr_mem_8_cns_douta_sho0),
      .shr_mem_8_cns_douta_sho1(shr_mem_8_cns_douta_sho1),
      .shr_mem_8_cns_S1_pff(shr_mem_8_cns_S1_iff),
      .din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_8_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_8_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_8_cns_S0_pff(shr_mem_8_cns_S0_iff)
    );
  double_buffeYeetf_9_cns_bctl double_buffeYeetf_9_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_9_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_9_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_9_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_9_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_9_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_9_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_9_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_9_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_9_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_9_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_9_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_9_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_9_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_9_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_9_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_9_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_9_cns_S0(shr_mem_9_cns_S0_dmo),
      .shr_mem_9_cns_R0(shr_mem_9_cns_R0),
      .shr_mem_9_cns_S1(shr_mem_9_cns_S1_dmo),
      .shr_mem_9_cns_R1(shr_mem_9_cns_R1),
      .shr_mem_9_cns_addra_shi0(shr_mem_9_cns_addra_shi0),
      .shr_mem_9_cns_addra_shi1(shr_mem_9_cns_addra_shi1),
      .shr_mem_9_cns_addrb_shi0(shr_mem_9_cns_addrb_shi0),
      .shr_mem_9_cns_addrb_shi1(shr_mem_9_cns_addrb_shi1),
      .shr_mem_9_cns_csa_n_shi0(shr_mem_9_cns_csa_n_shi0),
      .shr_mem_9_cns_csa_n_shi1(shr_mem_9_cns_csa_n_shi1),
      .shr_mem_9_cns_csb_n_shi0(shr_mem_9_cns_csb_n_shi0),
      .shr_mem_9_cns_csb_n_shi1(shr_mem_9_cns_csb_n_shi1),
      .shr_mem_9_cns_dinb_shi0(shr_mem_9_cns_dinb_shi0),
      .shr_mem_9_cns_dinb_shi1(shr_mem_9_cns_dinb_shi1),
      .shr_mem_9_cns_douta_sho0(shr_mem_9_cns_douta_sho0),
      .shr_mem_9_cns_douta_sho1(shr_mem_9_cns_douta_sho1),
      .shr_mem_9_cns_S1_pff(shr_mem_9_cns_S1_iff),
      .din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_9_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_9_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_9_cns_S0_pff(shr_mem_9_cns_S0_iff)
    );
  double_buffefnCNP10_cns_bctl double_buffefnCNP10_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_10_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_10_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_10_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_10_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_10_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_10_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_10_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_10_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_10_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_10_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_10_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_10_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_10_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_10_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_10_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_10_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_10_cns_S0(shr_mem_10_cns_S0_dmo),
      .shr_mem_10_cns_R0(shr_mem_10_cns_R0),
      .shr_mem_10_cns_S1(shr_mem_10_cns_S1_dmo),
      .shr_mem_10_cns_R1(shr_mem_10_cns_R1),
      .shr_mem_10_cns_addra_shi0(shr_mem_10_cns_addra_shi0),
      .shr_mem_10_cns_addra_shi1(shr_mem_10_cns_addra_shi1),
      .shr_mem_10_cns_addrb_shi0(shr_mem_10_cns_addrb_shi0),
      .shr_mem_10_cns_addrb_shi1(shr_mem_10_cns_addrb_shi1),
      .shr_mem_10_cns_csa_n_shi0(shr_mem_10_cns_csa_n_shi0),
      .shr_mem_10_cns_csa_n_shi1(shr_mem_10_cns_csa_n_shi1),
      .shr_mem_10_cns_csb_n_shi0(shr_mem_10_cns_csb_n_shi0),
      .shr_mem_10_cns_csb_n_shi1(shr_mem_10_cns_csb_n_shi1),
      .shr_mem_10_cns_dinb_shi0(shr_mem_10_cns_dinb_shi0),
      .shr_mem_10_cns_dinb_shi1(shr_mem_10_cns_dinb_shi1),
      .shr_mem_10_cns_douta_sho0(shr_mem_10_cns_douta_sho0),
      .shr_mem_10_cns_douta_sho1(shr_mem_10_cns_douta_sho1),
      .shr_mem_10_cns_S1_pff(shr_mem_10_cns_S1_iff),
      .din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_10_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_10_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_10_cns_S0_pff(shr_mem_10_cns_S0_iff)
    );
  double_buffefnCNP11_cns_bctl double_buffefnCNP11_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_11_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_11_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_11_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_11_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_11_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_11_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_11_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_11_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_11_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_11_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_11_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_11_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_11_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_11_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_11_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_11_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_11_cns_S0(shr_mem_11_cns_S0_dmo),
      .shr_mem_11_cns_R0(shr_mem_11_cns_R0),
      .shr_mem_11_cns_S1(shr_mem_11_cns_S1_dmo),
      .shr_mem_11_cns_R1(shr_mem_11_cns_R1),
      .shr_mem_11_cns_addra_shi0(shr_mem_11_cns_addra_shi0),
      .shr_mem_11_cns_addra_shi1(shr_mem_11_cns_addra_shi1),
      .shr_mem_11_cns_addrb_shi0(shr_mem_11_cns_addrb_shi0),
      .shr_mem_11_cns_addrb_shi1(shr_mem_11_cns_addrb_shi1),
      .shr_mem_11_cns_csa_n_shi0(shr_mem_11_cns_csa_n_shi0),
      .shr_mem_11_cns_csa_n_shi1(shr_mem_11_cns_csa_n_shi1),
      .shr_mem_11_cns_csb_n_shi0(shr_mem_11_cns_csb_n_shi0),
      .shr_mem_11_cns_csb_n_shi1(shr_mem_11_cns_csb_n_shi1),
      .shr_mem_11_cns_dinb_shi0(shr_mem_11_cns_dinb_shi0),
      .shr_mem_11_cns_dinb_shi1(shr_mem_11_cns_dinb_shi1),
      .shr_mem_11_cns_douta_sho0(shr_mem_11_cns_douta_sho0),
      .shr_mem_11_cns_douta_sho1(shr_mem_11_cns_douta_sho1),
      .shr_mem_11_cns_S1_pff(shr_mem_11_cns_S1_iff),
      .din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_11_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_11_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_11_cns_S0_pff(shr_mem_11_cns_S0_iff)
    );
  double_buffefnCNP12_cns_bctl double_buffefnCNP12_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_12_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_12_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_12_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_12_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_12_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_12_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_12_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_12_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_12_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_12_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_12_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_12_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_12_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_12_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_12_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_12_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_12_cns_S0(shr_mem_12_cns_S0_dmo),
      .shr_mem_12_cns_R0(shr_mem_12_cns_R0),
      .shr_mem_12_cns_S1(shr_mem_12_cns_S1_dmo),
      .shr_mem_12_cns_R1(shr_mem_12_cns_R1),
      .shr_mem_12_cns_addra_shi0(shr_mem_12_cns_addra_shi0),
      .shr_mem_12_cns_addra_shi1(shr_mem_12_cns_addra_shi1),
      .shr_mem_12_cns_addrb_shi0(shr_mem_12_cns_addrb_shi0),
      .shr_mem_12_cns_addrb_shi1(shr_mem_12_cns_addrb_shi1),
      .shr_mem_12_cns_csa_n_shi0(shr_mem_12_cns_csa_n_shi0),
      .shr_mem_12_cns_csa_n_shi1(shr_mem_12_cns_csa_n_shi1),
      .shr_mem_12_cns_csb_n_shi0(shr_mem_12_cns_csb_n_shi0),
      .shr_mem_12_cns_csb_n_shi1(shr_mem_12_cns_csb_n_shi1),
      .shr_mem_12_cns_dinb_shi0(shr_mem_12_cns_dinb_shi0),
      .shr_mem_12_cns_dinb_shi1(shr_mem_12_cns_dinb_shi1),
      .shr_mem_12_cns_douta_sho0(shr_mem_12_cns_douta_sho0),
      .shr_mem_12_cns_douta_sho1(shr_mem_12_cns_douta_sho1),
      .shr_mem_12_cns_S1_pff(shr_mem_12_cns_S1_iff),
      .din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_12_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_12_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_12_cns_S0_pff(shr_mem_12_cns_S0_iff)
    );
  double_buffefnCNP13_cns_bctl double_buffefnCNP13_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_13_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_13_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_13_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_13_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_13_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_13_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_13_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_13_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_13_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_13_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_13_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_13_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_13_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_13_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_13_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_13_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_13_cns_S0(shr_mem_13_cns_S0_dmo),
      .shr_mem_13_cns_R0(shr_mem_13_cns_R0),
      .shr_mem_13_cns_S1(shr_mem_13_cns_S1_dmo),
      .shr_mem_13_cns_R1(shr_mem_13_cns_R1),
      .shr_mem_13_cns_addra_shi0(shr_mem_13_cns_addra_shi0),
      .shr_mem_13_cns_addra_shi1(shr_mem_13_cns_addra_shi1),
      .shr_mem_13_cns_addrb_shi0(shr_mem_13_cns_addrb_shi0),
      .shr_mem_13_cns_addrb_shi1(shr_mem_13_cns_addrb_shi1),
      .shr_mem_13_cns_csa_n_shi0(shr_mem_13_cns_csa_n_shi0),
      .shr_mem_13_cns_csa_n_shi1(shr_mem_13_cns_csa_n_shi1),
      .shr_mem_13_cns_csb_n_shi0(shr_mem_13_cns_csb_n_shi0),
      .shr_mem_13_cns_csb_n_shi1(shr_mem_13_cns_csb_n_shi1),
      .shr_mem_13_cns_dinb_shi0(shr_mem_13_cns_dinb_shi0),
      .shr_mem_13_cns_dinb_shi1(shr_mem_13_cns_dinb_shi1),
      .shr_mem_13_cns_douta_sho0(shr_mem_13_cns_douta_sho0),
      .shr_mem_13_cns_douta_sho1(shr_mem_13_cns_douta_sho1),
      .shr_mem_13_cns_S1_pff(shr_mem_13_cns_S1_iff),
      .din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_13_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_13_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_13_cns_S0_pff(shr_mem_13_cns_S0_iff)
    );
  double_buffefnCNP14_cns_bctl double_buffefnCNP14_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_14_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_14_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_14_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_14_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_14_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_14_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_14_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_14_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_14_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_14_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_14_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_14_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_14_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_14_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_14_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_14_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_14_cns_S0(shr_mem_14_cns_S0_dmo),
      .shr_mem_14_cns_R0(shr_mem_14_cns_R0),
      .shr_mem_14_cns_S1(shr_mem_14_cns_S1_dmo),
      .shr_mem_14_cns_R1(shr_mem_14_cns_R1),
      .shr_mem_14_cns_addra_shi0(shr_mem_14_cns_addra_shi0),
      .shr_mem_14_cns_addra_shi1(shr_mem_14_cns_addra_shi1),
      .shr_mem_14_cns_addrb_shi0(shr_mem_14_cns_addrb_shi0),
      .shr_mem_14_cns_addrb_shi1(shr_mem_14_cns_addrb_shi1),
      .shr_mem_14_cns_csa_n_shi0(shr_mem_14_cns_csa_n_shi0),
      .shr_mem_14_cns_csa_n_shi1(shr_mem_14_cns_csa_n_shi1),
      .shr_mem_14_cns_csb_n_shi0(shr_mem_14_cns_csb_n_shi0),
      .shr_mem_14_cns_csb_n_shi1(shr_mem_14_cns_csb_n_shi1),
      .shr_mem_14_cns_dinb_shi0(shr_mem_14_cns_dinb_shi0),
      .shr_mem_14_cns_dinb_shi1(shr_mem_14_cns_dinb_shi1),
      .shr_mem_14_cns_douta_sho0(shr_mem_14_cns_douta_sho0),
      .shr_mem_14_cns_douta_sho1(shr_mem_14_cns_douta_sho1),
      .shr_mem_14_cns_S1_pff(shr_mem_14_cns_S1_iff),
      .din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_14_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_14_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_14_cns_S0_pff(shr_mem_14_cns_S0_iff)
    );
  double_buffefnCNP15_cns_bctl double_buffefnCNP15_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_addra_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .dout_15_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_15_rsc_addrb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_15_rsc_dinb_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_15_rsc_douta_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(dout_15_rsc_req_vz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_addra_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(8'b0),
      .din_15_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_15_rsc_addrb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_15_rsc_dinb_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_15_rsc_douta_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst(din_15_rsc_req_vz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst),
      .din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz(1'b0),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(dout_15_rsc_csa_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .dout_15_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(dout_15_rsc_rls_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud(din_15_rsc_csa_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud),
      .din_15_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud(din_15_rsc_rls_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_bud),
      .shr_mem_15_cns_S0(shr_mem_15_cns_S0_dmo),
      .shr_mem_15_cns_R0(shr_mem_15_cns_R0),
      .shr_mem_15_cns_S1(shr_mem_15_cns_S1_dmo),
      .shr_mem_15_cns_R1(shr_mem_15_cns_R1),
      .shr_mem_15_cns_addra_shi0(shr_mem_15_cns_addra_shi0),
      .shr_mem_15_cns_addra_shi1(shr_mem_15_cns_addra_shi1),
      .shr_mem_15_cns_addrb_shi0(shr_mem_15_cns_addrb_shi0),
      .shr_mem_15_cns_addrb_shi1(shr_mem_15_cns_addrb_shi1),
      .shr_mem_15_cns_csa_n_shi0(shr_mem_15_cns_csa_n_shi0),
      .shr_mem_15_cns_csa_n_shi1(shr_mem_15_cns_csa_n_shi1),
      .shr_mem_15_cns_csb_n_shi0(shr_mem_15_cns_csb_n_shi0),
      .shr_mem_15_cns_csb_n_shi1(shr_mem_15_cns_csb_n_shi1),
      .shr_mem_15_cns_dinb_shi0(shr_mem_15_cns_dinb_shi0),
      .shr_mem_15_cns_dinb_shi1(shr_mem_15_cns_dinb_shi1),
      .shr_mem_15_cns_douta_sho0(shr_mem_15_cns_douta_sho0),
      .shr_mem_15_cns_douta_sho1(shr_mem_15_cns_douta_sho1),
      .shr_mem_15_cns_S1_pff(shr_mem_15_cns_S1_iff),
      .din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(din_15_rsc_csb_n_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_pff(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_iff),
      .dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_pff(dout_15_rsc_csb_n_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst_buz_bud_iff),
      .shr_mem_15_cns_S0_pff(shr_mem_15_cns_S0_iff)
    );
  assign din_rsc_lz = din_rsc_lz_nWRITE_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_rsc_lz = dout_rsc_lz_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
  assign dout_rsc_z = dout_rsc_z_nREAD_BLOCK_OUTPUT_DTYPE_16_64_4_2_inst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    hls_target
// ------------------------------------------------------------------


module hls_target (
  clk, rst, input_rsc_z, input_rsc_vz, input_rsc_lz, weight_rsc_z, weight_rsc_vz,
      weight_rsc_lz, output_rsc_z, output_rsc_vz, output_rsc_lz, clamp_mem, scan_n,
      shift_n, slp_nret_n, slp_ret_n
);
  input clk;
  input rst;
  input [15:0] input_rsc_z;
  input input_rsc_vz;
  output input_rsc_lz;
  input [63:0] weight_rsc_z;
  input weight_rsc_vz;
  output weight_rsc_lz;
  output [1023:0] output_rsc_z;
  input output_rsc_vz;
  output output_rsc_lz;
  input clamp_mem;
  input scan_n;
  input shift_n;
  input slp_nret_n;
  input slp_ret_n;


  // Interconnect Declarations
  wire [511:0] dout_rsc_z_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst;
  wire dout_rsc_vz_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst;
  wire [63:0] dout_rsc_z_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst;
  wire dout_rsc_vz_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst;
  wire [511:0] input_rsc_z_nsystolic_array_inst;
  wire input_rsc_vz_nsystolic_array_inst;
  wire [63:0] weight_rsc_z_nsystolic_array_inst;
  wire weight_rsc_vz_nsystolic_array_inst;
  wire [1023:0] output_rsc_z_nsystolic_array_inst;
  wire output_rsc_vz_nsystolic_array_inst;
  wire [1023:0] din_rsc_z_ndouble_buffer_output_DTYPE_2_16_64_4_inst;
  wire din_rsc_vz_ndouble_buffer_output_DTYPE_2_16_64_4_inst;
  wire [1023:0] dout_rsc_z_ndouble_buffer_output_DTYPE_2_16_64_4_inst;
  wire din_rsc_lz_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst_bud;
  wire dout_rsc_lz_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst_bud;
  wire input_rsc_lz_nsystolic_array_inst_bud;
  wire din_rsc_lz_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst_bud;
  wire dout_rsc_lz_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst_bud;
  wire weight_rsc_lz_nsystolic_array_inst_bud;
  wire output_rsc_lz_nsystolic_array_inst_bud;
  wire din_rsc_lz_ndouble_buffer_output_DTYPE_2_16_64_4_inst_bud;
  wire dout_rsc_lz_ndouble_buffer_output_DTYPE_2_16_64_4_inst_bud;
  wire input_copy_unc_2;
  wire weight_copy_unc_2;
  wire output_copy_unc_2;


  // Interconnect Declarations for Component Instantiations 
  mgc_pipe_v10 #(.rscid(32'sd199),
  .width(32'sd512),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd1)) input_copy_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .ldin(input_rsc_lz_nsystolic_array_inst_bud),
      .vdin(input_rsc_vz_nsystolic_array_inst),
      .din(input_rsc_z_nsystolic_array_inst),
      .ldout(dout_rsc_lz_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst_bud),
      .vdout(dout_rsc_vz_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst),
      .dout(dout_rsc_z_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst),
      .sd(input_copy_unc_2)
    );
  mgc_pipe_v10 #(.rscid(32'sd200),
  .width(32'sd64),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd1)) weight_copy_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .ldin(weight_rsc_lz_nsystolic_array_inst_bud),
      .vdin(weight_rsc_vz_nsystolic_array_inst),
      .din(weight_rsc_z_nsystolic_array_inst),
      .ldout(dout_rsc_lz_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst_bud),
      .vdout(dout_rsc_vz_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst),
      .dout(dout_rsc_z_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst),
      .sd(weight_copy_unc_2)
    );
  mgc_pipe_v10 #(.rscid(32'sd201),
  .width(32'sd1024),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd1)) output_copy_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .ldin(din_rsc_lz_ndouble_buffer_output_DTYPE_2_16_64_4_inst_bud),
      .vdin(din_rsc_vz_ndouble_buffer_output_DTYPE_2_16_64_4_inst),
      .din(din_rsc_z_ndouble_buffer_output_DTYPE_2_16_64_4_inst),
      .ldout(output_rsc_lz_nsystolic_array_inst_bud),
      .vdout(output_rsc_vz_nsystolic_array_inst),
      .dout(output_rsc_z_nsystolic_array_inst),
      .sd(output_copy_unc_2)
    );
  double_buffer_input_DTYPE_64_16_4_1_3 double_buffer_input_DTYPE_64_16_4_1_3_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(input_rsc_z),
      .din_rsc_vz(input_rsc_vz),
      .din_rsc_lz(din_rsc_lz_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst_bud),
      .dout_rsc_z(dout_rsc_z_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst),
      .dout_rsc_vz(dout_rsc_vz_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst),
      .dout_rsc_lz(dout_rsc_lz_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst_bud),
      .clamp_mem(clamp_mem),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n)
    );
  double_buffer_weights_DTYPE_2_16_4_1_3 double_buffer_weights_DTYPE_2_16_4_1_3_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(weight_rsc_z),
      .din_rsc_vz(weight_rsc_vz),
      .din_rsc_lz(din_rsc_lz_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst_bud),
      .dout_rsc_z(dout_rsc_z_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst),
      .dout_rsc_vz(dout_rsc_vz_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst),
      .dout_rsc_lz(dout_rsc_lz_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst_bud),
      .clamp_mem(clamp_mem),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n)
    );
  systolic_array systolic_array_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_z(input_rsc_z_nsystolic_array_inst),
      .input_rsc_vz(input_rsc_vz_nsystolic_array_inst),
      .input_rsc_lz(input_rsc_lz_nsystolic_array_inst_bud),
      .weight_rsc_z(weight_rsc_z_nsystolic_array_inst),
      .weight_rsc_vz(weight_rsc_vz_nsystolic_array_inst),
      .weight_rsc_lz(weight_rsc_lz_nsystolic_array_inst_bud),
      .output_rsc_z(output_rsc_z_nsystolic_array_inst),
      .output_rsc_vz(output_rsc_vz_nsystolic_array_inst),
      .output_rsc_lz(output_rsc_lz_nsystolic_array_inst_bud)
    );
  double_buffer_output_DTYPE_2_16_64_4 double_buffer_output_DTYPE_2_16_64_4_inst
      (
      .clk(clk),
      .rst(rst),
      .din_rsc_z(din_rsc_z_ndouble_buffer_output_DTYPE_2_16_64_4_inst),
      .din_rsc_vz(din_rsc_vz_ndouble_buffer_output_DTYPE_2_16_64_4_inst),
      .din_rsc_lz(din_rsc_lz_ndouble_buffer_output_DTYPE_2_16_64_4_inst_bud),
      .dout_rsc_z(dout_rsc_z_ndouble_buffer_output_DTYPE_2_16_64_4_inst),
      .dout_rsc_vz(output_rsc_vz),
      .dout_rsc_lz(dout_rsc_lz_ndouble_buffer_output_DTYPE_2_16_64_4_inst_bud),
      .clamp_mem(clamp_mem),
      .scan_n(scan_n),
      .shift_n(shift_n),
      .slp_nret_n(slp_nret_n),
      .slp_ret_n(slp_ret_n)
    );
  assign input_rsc_lz = din_rsc_lz_ndouble_buffer_input_DTYPE_64_16_4_1_3_inst_bud;
  assign weight_rsc_lz = din_rsc_lz_ndouble_buffer_weights_DTYPE_2_16_4_1_3_inst_bud;
  assign output_rsc_lz = dout_rsc_lz_ndouble_buffer_output_DTYPE_2_16_64_4_inst_bud;
  assign output_rsc_z = dout_rsc_z_ndouble_buffer_output_DTYPE_2_16_64_4_inst;
endmodule



